--------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date:   15:30:00 05/20/2020
-- Design Name:
-- Module Name:   tms5220_tb.vhd
-- Project Name:  tms5220
-- Target Device:
-- Tool versions:
-- Description:
--
-- VHDL Test Bench Created by ISE for module: TMS5220
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes:
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation
-- simulation model.
--------------------------------------------------------------------------------
library ieee;
	use ieee.std_logic_1164.all;
	use ieee.std_logic_unsigned.all;
	use ieee.numeric_std.all;


entity tms5220_tb is
end tms5220_tb;

architecture behavior of tms5220_tb is
	--Inputs
	signal I_WSn    : std_logic := '0';
	signal I_RSn    : std_logic := '0';
	signal I_DATA   : std_logic := '0';
	signal I_TEST   : std_logic := '0';
	signal I_DBUS   : std_logic_vector(7 downto 0) := (others => '0');

	--Outputs
	signal CLK      : std_logic;
	signal O_RDYn   : std_logic;
	signal O_INTn   : std_logic;
	signal O_M0     : std_logic;
	signal O_M1     : std_logic;
	signal O_ADD8   : std_logic;
	signal O_ADD4   : std_logic;
	signal O_ADD2   : std_logic;
	signal O_ADD1   : std_logic;
	signal O_ROMCLK : std_logic;
	signal O_T11    : std_logic;
	signal O_IO     : std_logic;
	signal O_PRMOUT : std_logic;
	signal O_DBUS   : std_logic_vector(7 downto 0);
	signal O_SPKR   : signed(13 downto 0);

	signal
		current,
		index,
		offset,
		state        : integer := 0;

	constant MAXSOUNDS : integer := 141;
	type SIZE_ARRAY is array (0 to MAXSOUNDS-1) of integer;
	constant SIZES   : SIZE_ARRAY := (
		3651,248,141,117,138,133,150,89,120,72,147,112,154,47,415,456,375,402,153,221,157,128,182,124,325,217,182,182,497,356,288,407,335,486,
		351,398,201,217,173,194,123,104,244,178,144,116,109,109,78,109,150,247,164,192,201,88,128,166,84,59,72,69,47,84,97,172,166,72,116,84,78,
		84,103,247,128,72,53,372,335,497,502,212,323,209,250,311,276,300,325,91,103,108,486,455,242,343,438,373,214,358,407,492,404,422,491,261,
		352,280,197,299,382,213,214,164,328,331,63,270,172,111,102,67,86,103,111,129,116,141,128,159,304,434,435,418,316,329,461,203,179,479,316
	);

	constant DATALEN    : integer := 35598;
	type DATA_ARRAY is array (0 to DATALEN) of std_logic_vector(7 downto 0);
	constant DATA   : DATA_ARRAY := (
		-- speech data follows, CES phrase plus all Gauntlet sounds ID 8, 81..220, total audio 2m:41s
		x"60",x"80",x"D2",x"11",x"DC",x"54",x"4D",x"52",x"4A",x"B2",x"11",x"53",x"DF",x"98",x"2D",x"2D",x"4E",x"8D",x"63",x"62",x"A7",x"34",x"69",x"76",x"B3",x"72",x"1A",x"D2",x"64",x"B0",x"2C",x"D2",x"59",x"48",x"B3",x"81",x"B6",x"4A",x"67",x"25",x"29",x"86",x"C3",x"3D",x"A6",x"B4",x"64",x"38",x"16",x"0F",x"AB",x"1D",x"80",x"35",x"B7",x"1D",x"B0",x"E7",x"8E",x"03",x"76",x"BF",x"71",x"C0",x"1E",x"D7",x"0E",x"58",x"65",x"AB",x"48",x"5D",x"31",x"5B",x"75",x"EC",x"94",x"15",x"4E",x"35",x"6D",x"54",x"42",x"5A",x"04",x"4E",x"17",x"2B",x"0D",x"62",x"14",x"D2",x"9D",x"EC",x"38",x"C8",x"4E",x"65",x"79",x"9A",x"6A",x"A7",x"70",x"93",x"E5",x"E9",x"8E",x"95",x"CE",x"4C",x"8E",x"35",x"BB",x"4E",x"C6",x"54",x"8E",x"62",x"6E",x"CF",x"00",x"3F",x"BA",x"39",x"E0",x"6A",x"CB",x"B2",x"77",x"9B",x"E1",x"A6",x"94",x"8C",x"9B",x"58",x"58",x"9A",x"26",x"56",x"BE",x"CC",x"ED",x"CE",x"5A",x"C7",x"04",x"66",x"7A",x"19",x"44",x"1B",x"17",x"DA",x"65",x"5A",x"58",x"75",x"42",x"E4",x"BB",x"D8",x"72",x"CE",x"09",x"71",x"68",x"14",x"6B",x"D1",x"38",x"C5",x"B1",x"91",x"AF",x"65",x"92",x"90",x"C4",x"CA",x"F2",x"1E",x"71",x"42",x"9A",x"1A",x"E9",x"49",x"36",x"0A",x"69",x"99",x"A4",x"4B",x"39",x"55",x"ED",x"B9",x"61",x"B6",x"F6",x"12",x"24",x"A4",x"24",x"3E",x"51",x"DD",x"C8",x"35",x"92",x"67",x"9A",x"A5",x"45",x"D7",x"2C",x"91",x"AB",x"92",x"04",x"D0",x"D1",x"7C",x"B8",x"6A",x"D8",x"0E",x"F1",x"08",x"5A",x"2E",x"ED",x"78",x"14",x"35",x"98",x"9A",x"8E",x"AD",x"52",x"54",x"27",x"2A",x"B2",x"0A",x"5D",x"11",x"05",x"65",x"F9",x"B2",x"72",x"79",x"10",x"94",x"1D",x"CB",x"3A",x"E4",x"49",x"93",x"5B",x"8F",x"A3",x"91",x"B6",x"AA",x"8A",x"D5",x"2E",x"56",x"DC",x"B3",x"3A",x"4D",x"D9",x"5C",x"61",x"F5",x"16",x"3A",x"61",x"F9",x"04",x"35",x"5A",x"E8",x"84",x"9C",x"15",x"54",x"EB",x"29",x"55",x"56",x"5A",x"5C",x"B4",x"B7",x"84",x"DB",x"29",x"79",x"B2",x"65",x"11",x"1C",x"27",x"55",x"D1",x"B6",x"45",x"60",x"DD",x"D4",x"C4",x"10",x"11",x"22",x"F1",x"42",x"1B",x"83",x"87",x"51",x"24",x"31",x"7D",x"30",x"A9",x"C1",x"1D",x"45",x"0C",x"09",x"9B",x"65",x"78",x"1C",x"04",x"1C",x"13",x"22",x"80",x"EB",x"CB",x"19",x"F0",x"5C",x"86",x"00",x"BE",x"8F",x"50",x"C0",x"33",x"95",x"02",x"F8",x"7A",x"12",x"01",x"5F",x"A7",x"13",x"E0",x"B8",x"2D",x"00",x"E4",x"0E",x"47",x"62",x"D9",x"B6",x"5D",x"31",x"02",x"8A",x"CC",x"98",x"4A",x"45",x"F7",x"A8",x"3A",x"43",x"A9",x"94",x"23",x"92",x"72",x"AE",x"C5",x"56",x"8E",x"28",x"42",x"71",x"96",x"4A",x"D9",x"A2",x"B0",x"FA",x"C6",x"0A",x"55",x"B6",x"AC",x"56",x"2B",x"C9",x"54",x"56",x"73",x"47",x"05",x"2D",x"55",x"49",x"23",x"1B",x"6D",x"8C",x"58",x"43",x"9C",x"4D",x"47",x"D0",x"11",x"C0",x"8A",x"E9",x"A5",x"EE",x"DA",x"44",x"38",x"5A",x"97",x"7A",x"A8",x"62",x"45",x"5B",x"2C",x"80",x"1F",x"B2",x"04",x"F0",x"6B",x"85",x"00",x"7E",x"49",x"17",x"C0",x"2F",x"91",x"2D",x"AA",x"32",x"2C",x"B9",x"23",x"8D",x"A8",x"19",x"29",x"D7",x"8E",x"DC",x"E2",x"62",x"B4",x"DC",x"32",x"AA",x"8B",x"93",x"C1",x"76",x"F7",x"B8",x"2A",x"F6",x"9A",x"AA",x"22",x"ED",x"B0",x"D8",x"4B",x"8F",x"50",x"8F",x"ED",x"92",x"50",x"54",x"33",x"BD",x"75",x"48",x"63",x"66",x"3B",x"B3",x"BA",x"29",x"CF",x"45",x"68",x"53",x"16",x"95",x"22",x"67",x"96",x"0D",x"5D",x"54",x"CA",x"14",x"D8",x"2E",x"B5",x"76",x"A8",x"A3",x"E7",x"98",x"B0",x"B8",x"A2",x"CB",x"C6",x"C4",x"D4",x"E2",x"88",x"B6",x"38",x"75",x"77",x"95",x"A3",x"EA",x"28",x"D4",x"C2",x"DD",x"69",x"28",x"93",x"34",x"09",x"EF",x"5A",x"AD",x"AC",x"D9",x"D8",x"75",x"1D",x"B5",x"B2",x"16",x"71",x"CE",x"76",x"D8",x"CA",x"5E",x"C4",x"38",x"C7",x"45",x"29",x"7B",x"25",x"95",x"5C",x"87",x"A1",x"1A",x"8D",x"98",x"FD",x"55",x"98",x"66",x"44",x"63",x"96",x"B4",x"9A",x"9E",x"D9",x"2A",x"4C",x"32",x"32",x"03",x"D6",x"DA",x"60",x"C0",x"6E",x"A9",x"A1",x"1C",x"09",x"45",x"6F",x"44",x"85",x"6A",x"44",x"34",x"B9",x"A2",x"69",x"9A",x"28",x"D8",x"C7",x"1B",x"29",x"6B",x"A5",x"94",x"F3",x"34",x"CE",x"A1",x"9F",x"CE",x"55",x"55",x"6D",x"33",x"E0",x"96",x"28",x"01",x"BC",x"E1",x"29",x"80",x"E7",x"2B",x"19",x"B0",x"75",x"7A",x"2A",x"8B",x"91",x"92",x"58",x"47",x"A9",x"CA",x"9A",x"27",x"BC",x"6C",x"9B",x"26",x"6B",x"AE",x"94",x"8C",x"A2",x"BA",x"62",x"D8",x"CD",x"CC",x"89",x"6B",x"93",x"E4",x"CA",x"F4",x"D0",x"AE",x"8D",x"42",x"32",x"C2",x"A2",x"B8",x"2E",x"6B",x"E2",x"A8",x"B6",x"1C",x"BA",x"EE",x"51",x"A5",x"3B",x"85",x"E9",x"47",x"02",x"D1",x"6D",x"07",x"66",x"98",x"19",x"D1",x"6A",x"6D",x"99",x"61",x"36",x"62",x"EA",x"75",x"E4",x"C6",x"59",x"49",x"24",x"C7",x"96",x"9B",x"66",x"67",x"A5",x"AE",x"58",x"61",x"99",x"5D",x"0C",x"A7",x"12",x"A6",x"7D",x"0E",x"35",x"EA",x"4C",x"14",x"CE",x"39",x"D5",x"B1",x"B3",x"71",x"38",x"E7",x"CD",x"40",x"CB",x"26",x"66",x"5C",x"37",x"1C",x"AC",x"E2",x"98",x"61",x"2E",x"37",x"F4",x"8A",x"C3",x"AE",x"F9",x"66",x"9A",x"2C",x"09",x"5A",x"E6",x"A9",x"32",x"74",x"29",x"04",x"D8",x"EE",x"5A",x"00",x"DB",x"AC",x"11",x"60",x"D9",x"35",x"F5",x"0F",x"D3",x"CC",x"A4",x"A1",x"49",x"DB",x"6D",x"30",x"63",x"84",x"06",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"D7",x"CD",x"61",x"85",x"15",x"89",x"46",x"DE",x"03",x"97",x"54",x"3B",x"68",x"C5",x"08",x"54",x"1A",x"E5",x"C0",x"94",x"49",x"52",x"49",x"A6",x"22",x"57",x"06",x"25",x"19",x"D1",x"B2",x"5A",x"D1",x"A2",x"18",x"FB",x"AA",x"18",x"45",x"1F",x"62",x"92",x"E3",x"62",x"14",x"7D",x"B0",x"4A",x"8F",x"83",x"51",x"8C",x"26",x"C6",x"5B",x"31",x"46",x"3E",x"2A",x"87",x"6E",x"56",x"1C",x"79",x"8B",x"DC",x"B6",x"65",x"73",x"24",x"D5",x"EB",x"D8",x"46",x"AC",x"15",x"95",x"A8",x"ED",x"5D",x"B2",x"47",x"D0",x"12",x"57",x"64",x"CB",x"0A",x"FE",x"48",x"69",x"66",x"6E",x"6B",x"5C",x"B3",x"6D",x"45",x"A8",x"13",x"03",x"AC",x"7A",x"63",x"80",x"55",x"6F",x"0C",x"B0",x"DA",x"75",x"33",x"A7",x"35",x"73",x"D7",x"C6",x"CD",x"2E",x"C6",x"5B",x"35",x"3C",x"27",x"27",x"DA",x"69",x"D2",x"4E",x"5D",x"DC",x"24",x"BA",x"D8",x"DB",x"75",x"F3",x"2B",x"B3",x"B4",x"68",x"D7",x"25",x"EC",x"9A",x"55",x"72",x"63",x"99",x"B8",x"70",x"36",x"8F",x"B4",x"43",x"52",x"CF",x"C4",x"B2",x"DA",x"8E",x"4B",x"9B",x"45",x"B5",x"A8",x"36",x"29",x"1B",x"91",x"58",x"6A",x"53",x"BB",x"7C",x"16",x"24",x"EE",x"4D",x"49",x"F2",x"99",x"80",x"35",x"2A",x"31",x"01",x"76",x"CB",x"4E",x"D9",x"CA",x"C2",x"98",x"15",x"BB",x"65",x"63",x"08",x"73",x"6D",x"C2",x"91",x"8F",x"65",x"86",x"3E",x"2E",x"46",x"3E",x"9A",x"3A",x"56",x"25",x"68",x"C5",x"A8",x"1C",x"D4",x"19",x"A3",x"14",x"A3",x"50",x"62",x"B5",x"0B",x"57",x"56",x"0D",x"19",x"D1",x"0E",x"53",x"39",x"03",x"2B",x"BB",x"C7",x"36",x"C0",x"E9",x"33",x"0E",x"D8",x"E5",x"C6",x"01",x"AB",x"DD",x"38",x"60",x"8D",x"1B",x"07",x"AC",x"7E",x"63",x"80",x"35",x"AE",x"9B",x"DF",x"A3",x"32",x"7B",x"D7",x"1E",x"7E",x"0B",x"62",x"32",x"9D",x"A8",x"05",x"45",x"4B",x"44",x"96",x"5D",x"15",x"F5",x"A0",x"AA",x"EA",x"72",x"90",x"3B",x"63",x"9B",x"9A",x"A7",x"66",x"C3",x"8A",x"15",x"A1",x"66",x"3B",x"E5",x"CD",x"A9",x"4A",x"54",x"EC",x"52",x"8D",x"24",x"46",x"DD",x"09",x"D3",x"38",x"8A",x"98",x"54",x"C7",x"0A",x"CB",x"48",x"EC",x"3C",x"2E",x"45",x"AD",x"4D",x"51",x"6B",x"B1",x"63",x"B5",x"36",x"43",x"AD",x"21",x"4E",x"C4",x"52",x"15",x"0D",x"17",x"A7",x"62",x"4B",x"92",x"32",x"58",x"D2",x"48",x"CC",x"45",x"51",x"73",x"73",x"2A",x"D6",x"57",x"41",x"C5",x"25",x"8E",x"48",x"57",x"B4",x"38",x"3A",x"B7",x"42",x"75",x"B7",x"96",x"E8",x"E4",x"08",x"8D",x"C3",x"7B",x"71",x"A8",x"23",x"F4",x"B7",x"D2",x"AD",x"6E",x"8A",x"01",x"00",x"4C",x"3E",x"1B",x"31",x"F7",x"D8",x"4A",x"C5",x"A8",x"28",x"BC",x"65",x"31",x"95",x"23",x"B3",x"C2",x"B5",x"C4",x"50",x"35",x"47",x"46",x"DB",x"0A",x"54",x"6D",x"15",x"B7",x"77",x"32",x"52",x"75",x"50",x"D4",x"36",x"C9",x"42",x"D5",x"5E",x"73",x"E9",x"B4",x"4A",x"57",x"07",x"C3",x"9E",x"D6",x"8A",x"4A",x"5D",x"A2",x"A4",x"64",x"CB",x"6C",x"75",x"0B",x"92",x"E6",x"23",x"B9",x"D5",x"BD",x"B0",x"53",x"B5",x"A4",x"52",x"F7",x"46",x"AA",x"39",x"96",x"52",x"3D",x"1A",x"AA",x"F6",x"DA",x"34",x"F5",x"28",x"A8",x"94",x"EB",x"42",x"AC",x"B3",x"B4",x"B2",x"AB",x"ED",x"32",x"AD",x"76",x"A5",x"AA",x"96",x"04",x"B0",x"67",x"27",x"03",x"CE",x"4A",x"0B",x"E5",x"70",x"C8",x"31",x"4B",x"3A",x"54",x"23",x"A1",x"E8",x"0E",x"25",x"D7",x"14",x"85",x"D1",x"5D",x"88",x"54",x"A3",x"94",x"4C",x"84",x"69",x"36",x"6D",x"E0",x"EA",x"5D",x"E9",x"98",x"01",x"2B",x"94",x"0B",x"E0",x"A5",x"30",x"05",x"FC",x"9C",x"A1",x"80",x"5F",x"32",x"14",x"70",x"73",x"66",x"C9",x"8B",x"D4",x"48",x"9D",x"48",x"A5",x"88",x"DA",x"63",x"7C",x"2C",x"87",x"2A",x"A9",x"88",x"D6",x"B2",x"24",x"DA",x"2C",x"C5",x"DD",x"2C",x"B6",x"69",x"8B",x"64",x"4F",x"F5",x"A8",x"AE",x"49",x"52",x"A2",x"BC",x"02",x"AB",x"C6",x"48",x"AD",x"F2",x"92",x"ED",x"DA",x"22",x"31",x"B2",x"8A",x"92",x"EB",x"BA",x"41",x"8B",x"69",x"48",x"AE",x"1F",x"0E",x"55",x"B7",x"69",x"9A",x"A1",x"7B",x"54",x"9B",x"A2",x"25",x"C6",x"28",x"29",x"33",x"92",x"95",x"1A",x"A3",x"E4",x"4C",x"0D",x"27",x"61",x"A8",x"51",x"8D",x"B5",x"62",x"A5",x"A1",x"26",x"77",x"89",x"96",x"95",x"C6",x"12",x"32",x"25",x"4A",x"56",x"98",x"8A",x"CD",x"D2",x"48",x"25",x"61",x"29",x"2E",x"93",x"33",x"15",x"BB",x"AD",x"F8",x"48",x"C9",x"52",x"1C",x"8E",x"1E",x"BD",x"29",x"CA",x"76",x"B8",x"47",x"B1",x"16",x"AD",x"D8",x"66",x"EF",x"BB",x"56",x"43",x"53",x"BB",x"61",x"4C",x"6F",x"D2",x"72",x"25",x"D6",x"5E",x"D4",x"9C",x"CA",x"36",x"DA",x"5A",x"20",x"37",x"1E",x"C7",x"A4",x"EC",x"55",x"8B",x"35",x"34",x"8B",x"AC",x"D7",x"CC",x"50",x"95",x"CB",x"C6",x"51",x"D2",x"4C",x"2D",x"32",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"B0",x"BF",x"5B",x"15",x"63",x"77",x"9C",x"8A",x"EC",x"D4",x"D4",x"26",x"B6",x"02",x"AA",x"92",x"50",x"C0",x"8A",x"21",x"0A",x"58",x"A9",x"43",x"01",x"33",x"A6",x"A5",x"21",x"55",x"D3",x"08",x"4F",x"53",x"DC",x"52",x"5D",x"3C",x"3C",x"69",x"B3",x"6B",x"49",x"51",x"8B",x"BA",x"C3",x"2A",x"CE",x"59",x"23",x"E3",x"38",x"E0",x"EB",x"52",x"05",x"FC",x"B8",x"A1",x"80",x"9F",x"DB",x"18",x"F0",x"7D",x"79",x"1A",x"66",x"E8",x"0C",x"31",x"87",x"AD",x"1D",x"DE",x"34",x"28",x"6C",x"1E",x"AB",x"3A",x"4B",x"F5",x"B1",x"B5",x"EC",x"1A",x"22",x"A9",x"47",x"F2",x"70",x"4A",x"0A",x"97",x"58",x"29",x"C9",x"4D",x"DA",x"92",x"B5",x"1D",x"3B",x"37",x"0A",x"6E",x"CD",x"D0",x"E0",x"BC",x"C0",x"B5",x"CD",x"53",x"51",x"F2",x"0B",x"97",x"F2",x"68",x"4B",x"2D",x"A8",x"92",x"2B",x"AB",x"23",x"B5",x"28",x"2B",x"EE",x"8E",x"8C",x"1A",x"62",x"1F",x"3D",x"5C",x"62",x"8E",x"49",x"4C",x"0F",x"33",x"F6",x"2C",x"26",x"B1",x"5B",x"35",x"A4",x"D2",x"84",x"D8",x"2F",x"E6",x"B5",x"68",x"9A",x"92",x"98",x"C5",x"CE",x"B5",x"69",x"49",x"73",x"26",x"DF",x"F0",x"46",x"2D",x"CD",x"89",x"BD",x"23",x"52",x"95",x"24",x"05",x"89",x"0A",x"73",x"13",x"92",x"E2",x"DC",x"4D",x"D5",x"49",x"88",x"67",x"AA",x"4C",x"37",x"D9",x"69",x"28",x"31",x"55",x"C5",x"E3",x"24",x"3F",x"1F",x"8A",x"64",x"9F",x"92",x"82",x"72",x"D1",x"52",x"BC",x"49",x"89",x"6A",x"73",x"65",x"F5",x"24",x"2D",x"9D",x"7D",x"BB",x"D2",x"2C",x"2B",x"60",x"AC",x"6D",x"05",x"8C",x"B9",x"A3",x"80",x"B9",x"6E",x"0C",x"30",x"D7",x"CD",x"B8",x"67",x"BF",x"AE",x"49",x"CB",x"23",x"AA",x"5E",x"CD",x"BC",x"9A",x"8C",x"A8",x"68",x"0B",x"F7",x"9C",x"D2",x"E2",x"AC",x"B3",x"54",x"A2",x"4A",x"89",x"A3",x"DE",x"E0",x"90",x"A6",x"29",x"F6",x"AE",x"22",x"8C",x"EB",x"A6",x"38",x"A9",x"28",x"49",x"6E",x"1B",x"E2",x"24",x"34",x"BC",x"D5",x"55",x"49",x"8A",x"C8",x"E0",x"CC",x"24",x"25",x"2F",x"AA",x"93",x"2C",x"A3",x"96",x"B2",x"C8",x"18",x"B1",x"0C",x"93",x"AA",x"22",x"72",x"4D",x"23",x"68",x"AA",x"93",x"EE",x"16",x"8D",x"28",x"A9",x"89",x"6E",x"5A",x"35",x"AC",x"A4",x"2E",x"85",x"2E",x"8E",x"B6",x"92",x"FA",x"14",x"AB",x"29",x"DB",x"72",x"EA",x"53",x"CC",x"E6",x"98",x"C8",x"A9",x"CF",x"2E",x"46",x"75",x"62",x"A7",x"BF",x"49",x"D3",x"50",x"B6",x"14",x"DE",x"69",x"42",x"4D",x"D4",x"B2",x"4B",x"66",x"48",x"73",x"33",x"4B",x"61",x"9A",x"71",x"22",x"CC",x"6D",x"31",x"60",x"E5",x"0A",x"06",x"2C",x"D7",x"E1",x"D6",x"69",x"D3",x"5D",x"C5",x"0C",x"19",x"1B",x"75",x"8B",x"D0",x"A8",x"A8",x"0D",x"BA",x"32",x"4C",x"9D",x"01",x"F2",x"9B",x"30",x"33",x"77",x"A7",x"A8",x"64",x"A9",x"2A",x"94",x"55",x"8B",x"5A",x"D4",x"C8",x"20",x"73",x"A4",x"2A",x"13",x"3B",x"99",x"22",x"59",x"AA",x"A2",x"CA",x"4E",x"D6",x"BA",x"AD",x"2A",x"CA",x"32",x"34",x"AF",x"B4",x"BA",x"18",x"4B",x"B7",x"99",x"DC",x"EA",x"6C",x"CD",x"3D",x"A7",x"52",x"69",x"8A",x"53",x"B7",x"9C",x"9A",x"A5",x"29",x"5A",x"5D",x"EC",x"62",x"A7",x"A6",x"48",x"09",x"D7",x"8D",x"14",x"9A",x"86",x"43",x"42",x"73",x"91",x"00",x"9E",x"0E",x"13",x"C0",x"8F",x"A9",x"0C",x"F8",x"21",x"DD",x"F4",x"5D",x"B9",x"06",x"F6",x"E2",x"14",x"0C",x"BB",x"D9",x"24",x"B5",x"43",x"DE",x"A3",x"39",x"65",x"27",x"2E",x"45",x"CD",x"E2",x"5A",x"9D",x"B0",x"95",x"25",x"89",x"A7",x"6F",x"CA",x"52",x"D6",x"28",x"29",x"3A",x"1E",x"55",x"D3",x"92",x"BA",x"71",x"A8",x"42",x"45",x"AB",x"11",x"C1",x"E9",x"D5",x"14",x"33",x"65",x"94",x"B9",x"9D",x"52",x"36",x"C9",x"DE",x"56",x"51",x"52",x"95",x"58",x"54",x"BB",x"C6",x"15",x"4D",x"10",x"31",x"CE",x"6A",x"57",x"F4",x"D5",x"90",x"85",x"6B",x"1C",x"56",x"7B",x"AD",x"1D",x"6E",x"76",x"4C",x"61",x"62",x"B6",x"09",x"2B",x"49",x"79",x"D4",x"E9",x"A9",x"5C",x"B5",x"A5",x"35",x"88",x"AB",x"54",x"B5",x"12",x"B7",x"C8",x"49",x"39",x"A9",x"5D",x"5C",x"35",x"86",x"A7",x"C7",x"4A",x"F1",x"7C",x"9D",x"6A",x"6A",x"C5",x"00",x"AB",x"6D",x"A7",x"7F",x"A6",x"49",x"2F",x"89",x"93",x"82",x"12",x"4C",x"D4",x"23",x"4E",x"8A",x"52",x"61",x"9E",x"F0",x"24",x"21",x"89",x"85",x"F9",x"52",x"9B",x"86",x"2C",x"35",x"E2",x"35",x"6F",x"EA",x"F2",x"54",x"15",x"D6",x"B5",x"AE",x"28",x"73",x"73",x"68",x"B6",x"A4",x"A8",x"A9",x"A1",x"3D",x"58",x"1C",x"A5",x"BA",x"D5",x"89",x"F2",x"74",x"9C",x"DE",x"9E",x"D6",x"43",x"4C",x"56",x"4A",x"7A",x"4C",x"31",x"B2",x"3A",x"25",x"AF",x"46",x"25",x"A5",x"23",x"9B",x"32",x"4A",x"8E",x"92",x"65",x"6D",x"AA",x"2C",x"30",x"3B",x"CA",x"8A",x"00",x"4E",x"5C",x"17",x"C0",x"4F",x"19",x"02",x"F8",x"A1",x"4A",x"00",x"3F",x"67",x"29",x"E0",x"29",x"97",x"E2",x"57",x"25",x"9A",x"52",x"73",x"52",x"50",x"34",x"67",x"4A",x"55",x"35",x"41",x"76",x"10",x"EB",x"15",x"C6",x"84",x"39",x"40",x"8C",x"8D",x"65",x"13",x"05",x"2F",x"BE",x"EC",x"E1",x"43",x"1C",x"4A",x"D0",x"3A",x"4F",x"09",x"69",x"88",x"45",x"D3",x"54",x"BB",x"64",x"31",x"BA",x"6C",x"6B",x"AD",x"96",x"A7",x"20",x"3D",x"E6",x"71",x"5A",x"91",x"AC",x"77",x"8B",x"37",x"2D",x"45",x"D4",x"D9",x"4D",x"D1",x"24",x"14",x"51",x"76",x"25",x"66",x"BD",x"50",x"24",x"91",x"DD",x"94",x"51",x"5A",x"99",x"74",x"56",x"5A",x"C7",x"6E",x"65",x"B5",x"DC",x"E9",x"1D",x"BB",x"55",x"A3",x"1B",x"87",x"D9",x"EC",x"D0",x"8E",x"50",x"1D",x"45",x"96",x"D5",x"3D",x"43",x"4E",x"34",x"4B",x"0E",x"D3",x"AC",x"5E",x"D5",x"E6",x"A4",x"7D",x"23",x"4E",x"57",x"57",x"EC",x"F6",x"F5",x"30",x"D5",x"65",x"A2",x"D3",x"DF",x"42",x"55",x"98",x"39",x"29",x"69",x"CA",x"56",x"AE",x"51",x"65",x"64",x"C5",x"69",x"B7",x"79",x"DC",x"96",x"77",x"CB",x"13",x"11",x"96",x"5B",x"DE",x"83",x"34",x"77",x"C4",x"4A",x"79",x"F7",x"54",x"14",x"A5",x"B1",x"14",x"2D",x"6A",x"88",x"8C",x"AB",x"56",x"F6",x"CA",x"89",x"D5",x"1E",x"52",x"3D",x"16",x"05",x"4C",x"A5",x"10",x"40",x"CF",x"A4",x"0A",x"E8",x"AD",x"52",x"01",x"33",x"4F",x"1B",x"60",x"E5",x"59",x"03",x"CC",x"7E",x"6D",x"80",x"39",x"AE",x"0D",x"30",x"E7",x"8D",x"01",x"E6",x"B8",x"2E",x"65",x"B3",x"6A",x"EA",x"D1",x"B2",x"D4",x"C5",x"48",x"54",x"76",x"98",x"D2",x"65",x"6B",x"D1",x"91",x"71",x"52",x"9F",x"5C",x"44",x"6A",x"D4",x"09",x"7D",x"0C",x"19",x"6E",x"51",x"27",x"F4",x"D1",x"65",x"AB",x"E4",x"64",x"D7",x"27",x"93",x"6D",x"AC",x"93",x"54",x"1F",x"5D",x"0C",x"53",x"8E",x"36",x"7D",x"B4",x"39",x"46",x"72",x"5B",x"F5",x"3E",x"57",x"13",x"C5",x"15",x"D1",x"F8",x"54",x"4D",x"14",x"67",x"48",x"E3",x"CB",x"34",x"72",x"CC",x"25",x"BD",x"0B",x"3D",x"42",x"3E",x"87",x"35",x"AE",x"4F",x"30",x"DB",x"6D",x"D1",x"DA",x"DD",x"2A",x"62",x"B3",x"55",x"EB",x"7A",x"46",x"A0",x"CE",x"56",x"AD",x"DB",x"49",x"A5",x"BA",x"C8",x"74",x"A1",x"27",x"8D",x"F1",x"22",x"D3",x"85",x"1A",x"78",x"CE",x"93",x"5C",x"97",x"86",x"D2",x"86",x"34",x"72",x"5D",x"6E",x"86",x"D9",x"E2",x"D6",x"74",x"79",x"2A",x"C9",x"98",x"5D",x"F6",x"97",x"D2",x"81",x"E4",x"76",x"D0",x"DF",x"5C",x"A5",x"93",x"CA",x"01",x"00",x"00",x"40",x"7F",x"B3",x"E5",x"8A",x"39",x"07",x"01",x"4F",x"65",x"31",x"E0",x"87",x"4C",x"06",x"FC",x"98",x"29",x"80",x"9F",x"BA",x"04",x"F0",x"73",x"95",x"00",x"7E",x"AA",x"14",x"C0",x"0F",x"1D",x"02",x"38",x"32",x"24",x"25",x"23",x"11",x"8B",x"5F",x"EA",x"94",x"8E",x"8A",x"A4",x"B1",x"9D",x"43",x"36",x"2C",x"91",x"75",x"77",x"72",x"E9",x"70",x"48",x"71",x"93",x"08",x"01",x"6B",x"30",x"22",x"60",x"1D",x"42",x"04",x"AC",x"89",x"E4",x"8A",x"A1",x"90",x"6B",x"DB",x"91",x"2B",x"A7",x"43",x"F2",x"AB",x"58",x"A1",x"9C",x"0E",x"29",x"AE",x"6D",x"87",x"62",x"7A",x"24",x"9B",x"49",x"1C",x"8A",x"D9",x"90",x"F5",x"5A",x"B1",x"AB",x"E6",x"51",x"81",x"EE",x"C4",x"64",x"1A",x"95",x"54",x"77",x"1B",x"92",x"71",x"EE",x"1A",x"36",x"69",x"1B",x"DE",x"5E",x"25",x"64",x"A3",x"4E",x"6B",x"7A",x"E0",x"B4",x"AD",x"D8",x"AD",x"AE",x"4E",x"DA",x"37",x"63",x"B5",x"A6",x"78",x"ED",x"98",x"8C",x"5C",x"FA",x"1E",x"B4",x"74",x"A2",x"72",x"9B",x"5A",x"8A",x"E6",x"AA",x"26",x"69",x"6E",x"D1",x"9B",x"73",x"52",x"B9",x"B1",x"07",x"1B",x"B5",x"76",x"EC",x"FE",x"6E",x"D3",x"8A",x"3D",x"B6",x"00",x"8E",x"74",x"11",x"C0",x"0F",x"16",x"0C",x"F8",x"31",x"9C",x"01",x"BF",x"B8",x"31",x"E0",x"C7",x"4C",x"06",x"FC",x"12",x"C5",x"80",x"5F",x"A3",x"18",x"F0",x"4B",x"34",x"02",x"BE",x"A9",x"14",x"E6",x"54",x"5F",x"E5",x"1E",x"09",x"3D",x"3D",x"4C",x"A5",x"66",x"12",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"E4",x"8E",x"92",x"1D",x"92",x"59",x"42",x"DA",x"82",x"25",x"67",x"DB",x"6C",x"79",x"4F",x"D6",x"E8",x"99",x"B0",x"14",x"CD",x"72",x"B1",x"B5",x"C2",x"90",x"47",x"A5",x"AE",x"3A",x"2A",x"53",x"56",x"8C",x"3A",x"DB",x"31",x"6C",x"69",x"D7",x"92",x"AE",x"AB",x"60",x"A4",x"DD",x"6A",x"B8",x"8D",x"C3",x"95",x"F4",x"68",x"C5",x"3E",x"09",x"47",x"DC",x"A2",x"95",x"FA",x"26",x"49",x"4B",x"73",x"B2",x"EA",x"9D",x"54",x"F9",x"D1",x"46",x"B9",x"B9",x"55",x"95",x"D8",x"50",x"A5",x"6A",x"76",x"5D",x"EA",x"D2",x"14",x"71",x"C4",x"4D",x"59",x"52",x"DE",x"42",x"D5",x"A4",x"64",x"45",x"9B",x"3B",x"D7",x"DC",x"96",x"35",x"A5",x"EA",x"DC",x"F5",x"4A",x"DE",x"B4",x"8A",x"F1",x"36",x"0D",x"45",x"55",x"A6",x"42",x"33",x"D7",x"95",x"95",x"A6",x"88",x"D4",x"2C",x"06",x"6C",x"6A",x"C6",x"80",x"1F",x"3D",x"18",x"F0",x"7D",x"A7",x"71",x"A7",x"5C",x"27",x"8C",x"4C",x"46",x"1D",x"B1",x"33",x"34",x"C8",x"98",x"60",x"16",x"11",x"B2",x"4D",x"9C",x"D2",x"59",x"45",x"D0",x"2F",x"71",x"C9",x"BB",x"27",x"EA",x"18",x"B9",x"2D",x"9F",x"91",x"59",x"F5",x"64",x"B5",x"62",x"04",x"51",x"96",x"57",x"58",x"CA",x"EE",x"C5",x"58",x"4E",x"96",x"2B",x"A3",x"14",x"4F",x"5D",x"D5",x"A6",x"74",x"86",x"3B",x"BC",x"54",x"99",x"32",x"2A",x"2E",x"CD",x"88",x"19",x"B2",x"96",x"BC",x"49",x"AD",x"B5",x"30",x"4B",x"76",x"57",x"8F",x"A6",x"C8",x"AE",x"C1",x"C3",x"DD",x"E3",x"9A",x"24",x"0D",x"E1",x"35",x"5E",x"12",x"92",x"14",x"0B",x"66",x"A8",x"4E",x"4A",x"B2",x"1F",x"F0",x"95",x"D4",x"2D",x"4E",x"36",x"24",x"3B",x"12",x"8F",x"B8",x"4A",x"B1",x"8D",x"68",x"52",x"E2",x"8A",x"CD",x"2F",x"2C",x"AE",x"8B",x"13",x"C9",x"6A",x"71",x"BB",x"29",x"C9",x"34",x"32",x"DC",x"93",x"B4",x"AC",x"B2",x"50",x"8D",x"6A",x"D2",x"8A",x"61",x"94",x"DC",x"6A",x"4E",x"AA",x"47",x"66",x"12",x"B9",x"C6",x"A1",x"9D",x"5E",x"91",x"23",x"63",x"B1",x"69",x"5A",x"21",x"51",x"B7",x"2D",x"80",x"BD",x"A6",x"15",x"B0",x"E7",x"AD",x"02",x"D6",x"F8",x"6E",x"D1",x"EA",x"D7",x"19",x"22",x"B9",x"15",x"3D",x"3A",x"AA",x"65",x"E3",x"51",x"8E",x"CE",x"AA",x"B6",x"89",x"46",x"39",x"06",x"9B",x"F8",x"39",x"18",x"E5",x"E8",x"6C",x"92",x"6B",x"A3",x"15",x"A3",x"B0",x"49",x"B5",x"CD",x"92",x"F7",x"8C",x"2A",x"3D",x"32",x"42",x"9E",x"14",x"55",x"46",x"33",x"76",x"79",x"54",x"1C",x"E3",x"61",x"27",x"E5",x"4D",x"32",x"E6",x"96",x"95",x"54",x"36",x"4B",x"1C",x"E3",x"B5",x"53",x"95",x"8D",x"68",x"86",x"B5",x"76",x"8D",x"B7",x"E9",x"1D",x"9C",x"52",x"B5",x"36",x"85",x"37",x"F1",x"62",x"D3",x"85",x"E8",x"B6",x"CC",x"53",x"54",x"1F",x"B3",x"C8",x"19",x"DF",x"32",x"43",x"6E",x"AC",x"A7",x"3A",x"D9",x"8D",x"B9",x"B0",x"9C",x"C6",x"18",x"37",x"D6",x"2A",x"34",x"9A",x"63",x"DC",x"D8",x"06",x"AB",x"69",x"C7",x"0E",x"53",x"EF",x"A2",x"AC",x"53",x"DB",x"4D",x"BD",x"8B",x"A8",x"4E",x"AD",x"30",x"F5",x"A6",x"A2",x"52",x"B5",x"DD",x"D4",x"BC",x"9A",x"99",x"4F",x"55",x"73",x"35",x"6A",x"69",x"52",x"0B",x"2D",x"DD",x"29",x"89",x"98",x"6D",x"F6",x"77",x"EB",x"16",x"E1",x"72",x"CC",x"5D",x"BC",x"94",x"B9",x"38",x"71",x"75",x"96",x"98",x"6D",x"61",x"BB",x"34",x"45",x"AB",x"95",x"95",x"A5",x"D4",x"54",x"CB",x"19",x"5E",x"92",x"4B",x"DB",x"12",x"BB",x"E4",x"48",x"4A",x"4D",x"4F",x"64",x"52",x"2B",x"D3",x"35",x"CD",x"83",x"76",x"8D",x"28",x"D1",x"16",x"89",x"D6",x"D9",x"92",x"18",x"B0",x"EA",x"96",x"00",x"56",x"B9",x"60",x"C0",x"AE",x"1B",x"04",x"58",x"39",x"39",x"34",x"23",x"A1",x"EA",x"8C",x"28",x"D7",x"75",x"0B",x"E9",x"53",x"08",x"45",x"1F",x"24",x"75",x"7A",x"A2",x"52",x"43",x"10",x"12",x"E5",x"61",x"2B",x"F4",x"CB",x"85",x"A7",x"99",x"24",x"02",x"BC",x"A9",x"C9",x"80",x"9F",x"BD",x"18",x"F0",x"4B",x"A4",x"00",x"5E",x"C9",x"4C",x"79",x"A7",x"A6",x"6D",x"D9",x"B0",x"94",x"45",x"49",x"A5",x"6E",x"EC",x"50",x"65",x"AD",x"E5",x"36",x"B1",x"58",x"D7",x"A4",x"88",x"AB",x"39",x"36",x"6D",x"55",x"6A",x"6E",x"1E",x"C7",x"74",x"49",x"72",x"78",x"5B",x"4D",x"D3",x"27",x"49",x"11",x"95",x"A6",x"5C",x"5F",x"35",x"99",x"67",x"5B",x"32",x"43",x"53",x"60",x"DD",x"09",x"C7",x"8C",x"C3",x"21",x"7B",x"B5",x"64",x"37",x"F6",x"80",x"1C",x"D1",x"B2",x"D4",x"58",x"24",x"A5",x"6B",x"33",x"56",x"63",x"91",x"98",x"A9",x"A5",x"38",x"0C",x"D5",x"A9",x"3B",x"8F",x"E4",x"34",x"14",x"E3",x"69",x"56",x"B2",x"D3",x"50",x"6C",x"94",x"7A",x"C9",x"76",x"63",x"72",x"15",x"1A",x"AE",x"28",x"4C",x"C5",x"46",x"49",x"A4",x"15",x"B7",x"34",x"27",x"C5",x"15",x"91",x"CD",x"D6",x"B3",x"26",x"B5",x"97",x"71",x"DB",x"A8",x"92",x"94",x"19",x"D3",x"AD",x"3D",x"72",x"50",x"B7",x"43",x"31",x"77",x"4F",x"41",x"DE",x"0A",x"C9",x"98",x"35",x"87",x"EA",x"B2",x"24",x"7E",x"8B",x"11",x"0A",x"C9",x"99",x"D5",x"C3",x"95",x"1B",x"BB",x"1C",x"F6",x"0E",x"3F",x"6E",x"66",x"4E",x"FE",x"FF",
		x"60",x"0C",x"F8",x"21",x"9C",x"01",x"3F",x"A6",x"33",x"E0",x"A7",x"76",x"01",x"FC",x"D4",x"0C",x"06",x"E8",x"32",x"AC",x"EC",x"43",x"28",x"E4",x"76",x"AD",x"B2",x"4E",x"A6",x"90",x"3B",x"95",x"CA",x"3C",x"99",x"40",x"DD",x"46",x"6E",x"E3",x"14",x"02",x"B9",x"1B",x"B9",x"F5",x"93",x"09",x"D6",x"5E",x"A5",x"D2",x"4E",x"CA",x"D8",x"BD",x"91",x"42",x"DD",x"65",x"98",x"9B",x"D9",x"36",x"C0",x"AF",x"65",x"0A",x"78",x"7B",x"D3",x"00",x"6F",x"6E",x"0A",x"E0",x"B5",x"6D",x"06",x"DC",x"36",x"05",x"06",x"B8",x"D9",x"DD",x"00",x"EF",x"6C",x"19",x"E0",x"AD",x"EB",x"51",x"DE",x"B6",x"E1",x"02",x"B2",x"47",x"BE",x"1C",x"93",x"50",x"CC",x"1E",x"69",x"53",x"A2",x"91",x"53",x"69",x"C4",x"43",x"BA",x"B8",x"77",x"CD",x"16",x"36",x"11",x"9A",x"D6",x"95",x"9A",x"5F",x"79",x"6A",x"58",x"4E",x"1A",x"6E",x"96",x"E1",x"69",x"31",x"39",x"39",x"95",x"87",x"A5",x"66",x"6D",x"70",x"40",x"31",x"2E",x"0A",x"28",x"36",x"84",x"01",x"C5",x"95",x"00",x"80",x"03",x"8E",x"50",x"72",x"40",x"03",x"22",x"C3",x"CE",x"CA",x"2C",x"B2",x"60",x"0D",x"AB",x"EA",x"D0",x"8C",x"B5",x"B4",x"CC",x"A6",x"4A",x"D2",x"A7",x"D2",x"32",x"BA",x"6C",x"4D",x"EF",x"49",x"43",x"6F",x"72",x"24",x"AD",x"2B",x"35",x"2D",x"BB",x"F0",x"F0",x"15",x"9D",x"D4",x"A4",x"C3",x"C3",x"46",x"54",x"52",x"26",x"49",x"76",x"68",x"53",x"49",x"DE",x"50",x"C8",x"49",x"13",x"06",x"E9",x"BB",x"90",x"60",x"B1",x"19",x"C4",x"1F",x"CA",x"4A",x"D4",x"B1",x"11",x"7E",x"2A",x"35",x"16",x"3A",x"20",x"80",x"AB",x"D2",x"09",x"F0",x"55",x"E8",x"03",x"FF",
		x"60",x"AC",x"53",x"A2",x"AB",x"52",x"4D",x"B3",x"4E",x"A8",x"AE",x"74",x"B3",x"CC",x"5A",x"6E",x"BA",x"CA",x"CC",x"16",x"AB",x"99",x"DB",x"0C",x"35",x"DB",x"AA",x"60",x"B1",x"CB",x"D9",x"A3",x"98",x"84",x"E7",x"ED",x"24",x"9A",x"92",x"22",x"1B",x"DE",x"C9",x"6D",x"76",x"89",x"22",x"FF",x"C6",x"B0",x"85",x"2D",x"0A",x"E6",x"83",x"2A",x"6B",x"B7",x"38",x"9A",x"0B",x"89",x"A8",x"32",x"D2",x"A4",x"CF",x"24",x"A3",x"CA",x"28",x"92",x"1F",x"F1",x"8C",x"AA",x"A3",x"CE",x"B1",x"D9",x"BC",x"CA",x"8E",x"BE",x"A4",x"10",x"B6",x"89",x"12",x"86",x"AC",x"D8",x"59",x"27",x"8D",x"9B",x"B2",x"16",x"27",x"ED",x"BA",x"6E",x"CA",x"92",x"4D",x"B5",x"EB",x"BA",x"B9",x"68",x"56",x"91",x"6A",x"AA",x"D6",x"AC",x"59",x"45",x"AA",x"A9",x"DA",x"B2",x"71",x"14",x"8B",x"26",x"6A",x"2F",x"C9",x"C1",x"3A",x"CB",x"A2",x"93",x"67",x"C9",x"36",x"A2",x"FB",x"00",x"FF",
		x"60",x"02",x"68",x"41",x"8D",x"01",x"25",x"39",x"27",x"37",x"47",x"36",x"B6",x"58",x"92",x"BC",x"14",x"59",x"D5",x"F3",x"4D",x"F2",x"BC",x"35",x"8B",x"F2",x"3B",x"C9",x"B7",x"26",x"22",x"4A",x"E7",x"A4",x"D0",x"D8",x"F4",x"08",x"99",x"1D",x"12",x"9D",x"DD",x"DC",x"AB",x"A1",x"CB",x"54",x"D4",x"31",x"CE",x"45",x"21",x"E7",x"C5",x"D3",x"34",x"17",x"85",x"92",x"D7",x"32",x"B7",x"6C",x"ED",x"6A",x"91",x"22",x"9D",x"7D",x"AB",x"6B",x"85",x"6B",x"4F",x"D6",x"B6",x"6E",x"90",x"A6",x"23",x"45",x"D2",x"9A",x"49",x"BA",x"89",x"10",x"4D",x"6A",x"16",x"69",x"3B",x"43",x"24",x"A9",x"DA",x"94",x"1D",x"77",x"16",x"B7",x"EC",x"D0",x"66",x"D2",x"58",x"9D",x"92",x"9B",x"2C",x"63",x"8D",x"8A",x"F9",x"00",x"FF",
		x"60",x"04",x"48",x"C2",x"DC",x"A5",x"B1",x"92",x"BB",x"45",x"5A",x"13",x"85",x"81",x"56",x"A1",x"69",x"4C",x"18",x"3A",x"78",x"3B",x"67",x"09",x"41",x"6C",x"A8",x"35",x"DC",x"3A",x"84",x"79",x"A2",x"46",x"C8",x"A3",x"16",x"97",x"AC",x"24",x"ED",x"4D",x"5A",x"52",x"82",x"B0",x"6E",x"D6",x"6D",x"69",x"11",x"26",x"B6",x"55",x"65",x"64",x"4D",x"1B",x"73",x"F5",x"DC",x"91",x"0F",x"69",x"4C",x"35",x"73",x"5A",x"D9",x"85",x"32",x"F7",x"D4",x"69",x"D5",x"10",x"46",x"54",x"53",x"A7",x"35",x"93",x"2B",x"51",x"CD",x"E2",x"D6",x"4F",x"6E",x"44",x"35",x"4D",x"CA",x"B0",x"B8",x"12",x"D6",x"D4",x"4E",x"D3",x"92",x"46",x"98",x"33",x"3B",x"4D",x"93",x"2B",x"71",x"CD",x"EC",x"34",x"0F",x"AE",x"24",x"3D",x"93",x"DD",x"5A",x"99",x"92",x"CF",x"54",x"71",x"5B",x"15",x"4A",x"3E",x"5B",x"86",x"EC",x"56",x"71",x"56",x"3B",x"E9",x"07",x"FF",
		x"60",x"08",x"C8",x"D6",x"9C",x"02",x"2E",x"96",x"AB",x"52",x"B8",x"AA",x"86",x"48",x"F5",x"57",x"76",x"9B",x"9A",x"22",x"35",x"36",x"8C",x"AD",x"6A",x"8A",x"65",x"DF",x"74",x"D2",x"BA",x"29",x"51",x"69",x"2B",x"88",x"A7",x"A4",x"CC",x"FA",x"AD",x"24",x"9C",x"93",x"72",x"93",x"B7",x"82",x"68",x"76",x"29",x"74",x"9D",x"4A",x"92",x"25",x"A5",x"B4",x"B5",x"2B",x"50",x"57",x"97",x"DA",x"A7",x"AA",x"14",x"5A",x"55",x"5A",x"DF",x"23",x"52",x"74",x"55",x"E9",x"7D",x"37",x"2F",x"B5",x"55",x"65",x"08",x"43",x"AD",x"42",x"57",x"A6",x"31",x"76",x"8E",x"36",x"DD",x"98",x"A6",x"D4",x"B1",x"4A",x"6D",x"55",x"98",x"53",x"C7",x"2C",x"97",x"4D",x"61",x"4E",x"1D",x"2B",x"5D",x"36",x"B9",x"39",x"0D",x"AC",x"74",x"DD",x"E5",x"D6",x"34",x"B0",x"D2",x"AC",x"37",x"59",x"7D",x"C1",x"75",x"0D",x"93",x"0F",x"FF",
		x"60",x"08",x"C8",x"C6",x"9C",x"02",x"04",x"08",x"33",x"2C",x"65",x"61",x"A5",x"46",x"4E",x"94",x"96",x"C5",x"15",x"6E",x"D9",x"51",x"46",x"96",x"F2",x"98",x"7B",x"56",x"19",x"59",x"F6",x"EB",x"16",x"59",x"67",x"14",x"29",x"B6",x"BB",x"F7",x"94",x"51",x"A5",x"52",x"16",x"D9",x"53",x"47",x"93",x"4A",x"A9",x"47",x"57",x"1D",x"7D",x"1E",x"66",x"5E",x"13",x"65",x"0C",x"B9",x"B8",x"45",x"4D",x"99",x"31",x"E6",x"AA",x"61",x"3D",x"51",x"C6",x"98",x"93",x"7A",x"64",x"47",x"1D",x"63",x"89",x"6A",x"5E",x"5D",x"A5",x"4D",x"C5",x"A9",x"7B",x"F5",x"98",x"32",x"65",x"CF",x"56",x"53",x"65",x"DA",x"5C",x"8C",x"6A",x"F4",x"4C",x"69",x"4B",x"F1",x"4A",x"D1",x"B5",x"B8",x"2D",x"D5",x"AA",x"B8",x"C7",x"E3",x"B0",x"D6",x"20",x"EA",x"E2",x"4B",x"D0",x"8A",x"83",x"44",x"45",x"9A",x"02",x"B2",x"98",x"20",x"69",x"D9",x"A2",x"C8",x"6A",x"A3",x"36",x"67",x"10",x"41",x"AB",x"4F",x"68",x"E5",x"42",x"EA",x"01",x"FF",
		x"60",x"08",x"58",x"22",x"8D",x"00",x"47",x"55",x"10",x"E0",x"48",x"57",x"02",x"6C",x"DD",x"4E",x"80",x"29",x"53",x"4B",x"5C",x"BC",x"98",x"F8",x"D6",x"1D",x"71",x"31",x"C6",x"1E",x"3D",x"77",x"64",x"DD",x"87",x"A8",x"E6",x"93",x"51",x"76",x"1F",x"A2",x"96",x"4B",x"5A",x"DF",x"53",x"B0",x"B8",x"AF",x"31",x"47",x"5B",x"2C",x"E6",x"39",x"07",x"80",x"00",x"E5",x"50",x"10",x"60",x"A8",x"0B",x"02",x"2C",x"35",x"41",x"80",x"A3",x"32",x"08",x"B0",x"54",x"3B",x"01",x"96",x"28",x"47",x"C0",x"E6",x"EE",x"08",x"B8",x"2A",x"1D",x"1E",x"FF",
		x"60",x"08",x"98",x"26",x"8D",x"00",x"4B",x"86",x"12",x"60",x"89",x"D0",x"10",x"75",x"55",x"2C",x"5C",x"B5",x"4A",x"9C",x"A2",x"4A",x"4C",x"46",x"1D",x"71",x"C9",x"EE",x"E2",x"5D",x"67",x"C5",x"D5",x"95",x"B9",x"E6",x"9C",x"91",x"14",x"57",x"EA",x"9A",x"53",x"4A",x"9E",x"6D",x"AA",x"4B",x"5C",x"51",x"75",x"14",x"AE",x"61",x"51",x"29",x"95",x"39",x"B8",x"2A",x"C7",x"94",x"51",x"57",x"9B",x"EA",x"12",x"77",x"46",x"57",x"63",x"89",x"6A",x"2D",x"19",x"43",x"0B",x"E5",x"22",x"B1",x"38",x"4D",x"4D",x"86",x"B2",x"C9",x"1C",x"37",x"55",x"25",x"6A",x"EC",x"F3",x"DC",x"54",x"8D",x"AA",x"52",x"CC",x"37",x"4B",x"D1",x"AC",x"2A",x"55",x"4F",x"AD",x"D9",x"88",x"0A",x"57",x"3D",x"B5",x"25",x"2B",x"C2",x"52",x"4D",x"1F",x"FF",
		x"60",x"A9",x"28",x"5E",x"D4",x"AB",x"AB",x"8C",x"74",x"38",x"13",x"C9",x"5A",x"33",x"92",x"11",x"5C",x"D8",x"73",x"C9",x"48",x"BA",x"37",x"91",x"EC",x"25",x"23",x"E9",x"4E",x"59",x"7A",x"E6",x"8C",x"7C",x"18",x"16",x"9E",x"99",x"DD",x"9A",x"15",x"4C",x"C0",x"67",x"4D",x"19",x"56",x"0A",x"05",x"9A",x"D6",x"7A",x"00",x"00",x"06",x"4C",x"16",x"8A",x"80",x"61",x"59",x"10",x"D0",x"8C",x"29",x"02",x"B2",x"76",x"01",x"00",x"78",x"FF",
		x"60",x"6A",x"48",x"9C",x"B2",x"DC",x"6D",x"9B",x"D6",x"4B",x"2E",x"B3",x"8C",x"35",x"F2",x"16",x"3C",x"49",x"6C",x"F1",x"C8",x"4B",x"F1",x"24",x"CF",x"29",x"23",x"2B",x"A1",x"C2",x"25",x"C6",x"8E",x"34",x"DB",x"8D",x"50",x"9D",x"32",x"D2",x"EC",x"D6",x"34",x"A3",x"CA",x"48",x"B3",x"5B",x"D3",x"88",x"2A",x"23",x"CB",x"76",x"4D",x"23",x"AA",x"8C",x"2C",x"DB",x"35",x"CD",x"A8",x"32",x"F2",x"E2",x"D6",x"34",x"62",x"F2",x"A8",x"4A",x"6E",x"37",x"CD",x"B2",x"A3",x"69",x"A1",x"C2",x"D8",x"E7",x"8C",x"B6",x"87",x"70",x"35",x"5F",x"3C",x"FA",x"1E",x"52",x"C5",x"7C",x"C9",x"18",x"46",x"70",x"65",x"8B",x"45",x"63",x"1C",x"5E",x"45",x"22",x"66",x"B5",x"69",x"3A",x"65",x"09",x"5F",x"14",x"96",x"26",x"54",x"A4",x"BC",x"92",x"59",x"8A",x"22",x"0B",x"CB",x"32",x"66",x"C9",x"9A",x"5C",x"AD",x"E3",x"A8",x"35",x"2B",x"36",x"B5",x"AA",x"2D",x"D6",x"62",x"44",x"44",x"B2",x"F2",x"03",x"FF",
		x"60",x"0C",x"18",x"C2",x"8D",x"00",x"4B",x"B8",x"A6",x"A4",x"C7",x"14",x"95",x"A8",x"52",x"C2",x"62",x"C5",x"23",x"27",x"CA",x"08",x"6B",x"E2",x"90",x"6E",x"3B",x"2B",x"68",x"59",x"5D",x"AD",x"2B",x"AF",x"B0",x"65",x"57",x"D3",x"6E",x"BC",x"A2",x"96",x"43",x"4D",x"A6",x"CE",x"4A",x"6A",x"29",x"35",x"AE",x"3A",x"2B",x"AB",x"39",x"5D",x"A5",x"AA",x"AE",x"A2",x"46",x"57",x"D3",x"A9",x"32",x"EA",x"1A",x"8A",x"55",x"6A",x"4C",x"EB",x"9A",x"1D",x"62",x"F5",x"C9",x"A1",x"2F",x"D6",x"48",x"A8",x"AB",x"BA",x"A9",x"1A",x"15",x"85",x"AE",x"E6",x"A6",x"6A",x"44",x"15",x"BB",x"A9",x"9B",x"AB",x"32",x"36",x"8C",x"69",x"66",x"29",x"46",x"C5",x"28",x"E7",x"EA",x"E5",x"01",x"FF",
		x"60",x"04",x"60",x"26",x"83",x"01",x"46",x"99",x"84",x"7E",x"E8",x"10",x"25",x"CB",x"54",x"8A",x"6A",x"8D",x"55",x"A7",x"CE",x"48",x"9A",x"63",x"E3",x"E8",x"35",x"23",x"28",x"49",x"C4",x"2A",x"57",x"37",x"3F",x"55",x"F4",x"4C",x"5F",x"59",x"82",x"D8",x"B0",x"32",x"6C",x"53",x"48",x"C2",x"40",x"AF",x"B0",x"AC",x"21",x"F3",x"8D",x"B5",x"22",x"9C",x"B6",x"22",x"46",x"0B",x"CA",x"70",x"36",x"AA",x"90",x"25",x"C2",x"A3",x"E9",x"EA",x"A2",x"0B",x"AF",x"D0",x"59",x"AB",x"CF",x"2A",x"3D",x"93",x"57",x"AF",x"31",x"AB",x"8E",x"08",x"5E",x"35",x"A6",x"A8",x"C6",x"C3",x"65",x"D3",x"98",x"13",x"9F",x"F4",x"E0",x"4E",x"63",x"89",x"A2",x"33",x"9D",x"5B",x"97",x"25",x"8A",x"8E",x"34",x"5A",x"5D",x"D6",x"A0",x"2A",x"CA",x"79",x"51",x"59",x"83",x"9A",x"08",x"97",x"45",x"61",x"F3",x"76",x"22",x"54",x"57",x"87",x"C9",x"EB",x"4D",x"37",x"59",x"1D",x"76",x"6F",x"27",x"43",x"78",x"B3",x"59",x"BC",x"9D",x"0C",x"D1",x"2D",x"0F",x"FF",
		x"60",x"0B",x"E8",x"32",x"6C",x"03",x"1B",x"D8",x"C0",x"06",x"36",x"B0",x"81",x"0D",x"6C",x"60",x"03",x"1B",x"D8",x"C0",x"06",x"36",x"B0",x"81",x"0D",x"6C",x"60",x"03",x"1B",x"D8",x"C0",x"06",x"36",x"B0",x"81",x"0D",x"6C",x"60",x"03",x"1B",x"D8",x"C0",x"06",x"36",x"F0",x"00",x"FF",
		x"60",x"04",x"A8",x"45",x"82",x"01",x"B5",x"46",x"28",x"A0",x"94",x"70",x"06",x"A4",x"A2",x"11",x"34",x"7F",x"D5",x"79",x"24",x"55",x"D0",x"42",x"AB",x"A4",x"CD",x"58",x"C9",x"8C",x"33",x"4D",x"B2",x"A2",x"14",x"33",x"8E",x"52",x"ED",x"8C",x"5C",x"8C",x"B4",x"C2",x"34",x"B2",x"F1",x"30",x"53",x"0C",x"F5",x"CA",x"D8",x"CB",x"CA",x"D6",x"2D",x"3A",x"1A",x"2E",x"A7",x"38",x"95",x"28",x"8F",x"3C",x"FC",x"9A",x"55",x"2C",x"A3",x"F2",x"88",x"4A",x"10",x"F5",x"CC",x"D9",x"23",x"29",x"DE",x"4C",x"53",x"67",x"97",x"34",x"FB",x"70",x"75",x"4B",x"5D",x"B2",x"E2",x"D4",x"22",x"BC",x"62",x"CA",x"8B",x"37",x"F1",x"F4",x"5A",x"A9",x"AE",x"49",x"D4",x"C2",x"EB",x"86",x"A8",x"78",x"56",x"CF",x"5A",x"9C",x"D2",x"1A",x"D4",x"CC",x"6D",x"B1",x"EA",x"BD",x"53",x"B7",x"74",x"C5",x"08",x"F0",x"DA",x"02",x"01",x"C1",x"A9",x"13",x"20",x"7A",x"55",x"93",x"47",x"95",x"99",x"2E",x"91",x"42",x"E1",x"FB",x"98",x"78",x"CC",x"6C",x"45",x"0C",x"9D",x"6E",x"B2",x"A4",x"15",x"29",x"74",x"98",x"EA",x"EC",x"56",x"A4",x"D8",x"A6",x"E1",x"93",x"47",x"99",x"63",x"9A",x"86",x"CD",x"5E",x"55",x"F5",x"6E",x"9A",x"B6",x"7A",x"D4",x"2D",x"98",x"68",x"F8",x"EC",x"D1",x"74",x"69",x"62",x"AD",x"A5",x"52",x"9B",x"45",x"BA",x"05",x"C6",x"0E",x"5D",x"74",x"A1",x"2A",x"52",x"29",x"74",x"C9",x"9B",x"AA",x"59",x"A5",x"D4",x"17",x"6B",x"2A",x"AE",x"35",x"C3",x"D8",x"BC",x"88",x"86",x"57",x"0A",x"4E",x"F3",x"AE",x"2A",x"D4",x"A6",x"F5",x"C5",x"71",x"98",x"F4",x"E2",x"D6",x"27",x"27",x"E9",x"56",x"4B",x"DA",x"90",x"9C",x"45",x"8A",x"AC",x"4D",x"63",x"30",x"91",x"A9",x"94",x"D5",x"4C",x"DE",x"44",x"95",x"60",x"16",x"33",x"7A",x"5D",x"95",x"86",x"B6",x"DD",x"E0",x"AD",x"55",x"98",x"07",x"2E",x"43",x"B0",x"5E",x"ED",x"94",x"B8",x"0D",x"29",x"64",x"B8",x"D1",x"BA",x"31",x"95",x"6C",x"AE",x"AE",x"DD",x"C7",x"54",x"B3",x"AA",x"44",x"74",x"1B",x"73",x"4F",x"61",x"64",x"BE",x"76",x"CC",x"C3",x"BB",x"A1",x"F9",x"DA",x"31",x"CF",x"E0",x"86",x"EA",x"6B",x"C7",x"32",x"9C",x"19",x"85",x"57",x"1E",x"4B",x"0F",x"E6",x"14",x"DE",x"74",x"AC",x"2D",x"67",x"88",x"E9",x"B2",x"B1",x"D7",x"E0",x"A1",x"E5",x"4B",x"DB",x"56",x"A2",x"B7",x"86",x"2F",x"6D",x"53",x"89",x"D1",x"E1",x"BA",x"76",x"CC",x"C5",x"57",x"59",x"6A",x"D3",x"31",x"67",x"5F",x"65",x"A9",x"ED",x"C6",x"52",x"7C",x"54",x"06",x"B7",x"6D",x"4B",x"B1",x"56",x"95",x"DC",x"B4",x"AD",x"D9",x"79",x"A7",x"F1",x"D2",x"B2",x"27",x"1B",x"E5",x"8E",x"4B",x"DD",x"91",x"8C",x"67",x"B8",x"B4",x"01",x"20",x"40",x"E5",x"A5",x"08",x"98",x"2A",x"04",x"01",x"43",x"B8",x"3E",x"FF",
		x"60",x"6E",x"32",x"25",x"82",x"24",x"56",x"B7",x"31",x"D9",x"68",x"15",x"E9",x"3A",x"FA",x"6C",x"A2",x"9C",x"7C",x"ED",x"E8",x"8A",x"B0",x"1E",x"96",x"35",x"A3",x"4D",x"DC",x"E7",x"88",x"9B",x"96",x"36",x"73",x"DB",x"45",x"89",x"5B",x"BA",x"CA",x"64",x"1B",x"B5",x"8D",x"99",x"8B",x"E8",x"76",x"56",x"3B",x"40",x"00",x"1F",x"54",x"4A",x"95",x"BC",x"A9",x"7B",x"D5",x"1E",x"65",x"F4",x"16",x"66",x"D9",x"66",x"D4",x"51",x"55",x"B9",x"44",x"E3",x"51",x"47",x"33",x"2E",x"92",x"8B",x"4B",x"ED",x"C5",x"84",x"AB",x"C5",x"49",x"75",x"A0",x"E6",x"2D",x"19",x"27",x"54",x"56",x"58",x"A6",x"54",x"DC",x"50",x"6B",x"E1",x"99",x"D2",x"71",x"42",x"A5",x"A5",x"47",x"F1",x"D8",x"75",x"B9",x"D7",x"A6",x"A1",x"1B",x"27",x"E4",x"DE",x"BA",x"86",x"B6",x"AA",x"54",x"C6",x"54",x"26",x"92",x"8D",x"43",x"1D",x"4D",x"B9",x"4A",x"54",x"71",x"75",x"D0",x"69",x"E1",x"61",x"47",x"D5",x"51",x"AB",x"79",x"84",x"1C",x"51",x"45",x"61",x"6E",x"54",x"75",x"58",x"E5",x"B9",x"7B",x"68",x"D5",x"11",x"55",x"E0",x"E6",x"AE",x"D5",x"18",x"00",x"40",x"00",x"D5",x"2B",x"BB",x"BA",x"26",x"13",x"32",x"6D",x"9D",x"FA",x"68",x"D4",x"AC",x"62",x"56",x"1B",x"B3",x"16",x"57",x"CB",x"D5",x"66",x"CA",x"4A",x"4D",x"C4",x"5A",x"B7",x"B1",x"5A",x"73",x"41",x"6F",x"3B",x"BA",x"AA",x"CC",x"9C",x"63",x"F5",x"E8",x"9B",x"72",x"75",x"8A",x"2D",x"6A",x"4F",x"5C",x"DC",x"3D",x"6B",x"81",x"00",x"7A",x"10",x"17",x"40",x"8D",x"22",x"29",x"2D",x"35",x"DC",x"4C",x"2D",x"87",x"CC",x"57",x"8A",x"0A",x"F3",x"9A",x"B2",x"D0",x"30",x"C2",x"3D",x"6B",x"CB",x"53",x"25",x"77",x"AB",x"2E",x"A3",x"48",x"81",x"32",x"73",x"1A",x"8D",x"B2",x"66",x"16",x"AD",x"9A",x"3D",x"AA",x"EA",x"58",x"24",x"7B",x"C9",x"68",x"9A",x"13",x"21",x"EF",x"25",x"65",x"E8",x"CD",x"02",x"84",x"DB",x"18",x"60",x"54",x"51",x"03",x"8C",x"55",x"51",x"86",x"9C",x"58",x"2C",x"BC",x"4E",x"1A",x"52",x"03",x"AF",x"F0",x"56",x"6D",x"4E",x"9D",x"34",x"42",x"DA",x"B4",x"39",x"56",x"72",x"37",x"4F",x"DB",x"96",x"10",x"35",x"34",x"3C",x"69",x"59",x"93",x"D6",x"30",x"37",x"B9",x"69",x"2D",x"86",x"5C",x"C6",x"2D",x"9B",x"B5",x"1A",x"F4",x"74",x"89",x"D3",x"E6",x"6C",x"25",x"4D",x"22",x"76",x"99",x"42",x"D2",x"90",x"B2",x"AC",x"6D",x"0C",x"DE",x"83",x"D3",x"B6",x"8C",x"31",x"D8",x"48",x"09",x"EB",x"DA",x"E6",x"60",x"23",x"D4",x"B4",x"5B",x"59",x"82",x"89",x"74",x"95",x"ED",x"61",x"0B",x"35",x"82",x"C8",x"5B",x"BB",x"C3",x"DB",x"2C",x"15",x"4D",x"63",x"56",x"67",x"AB",x"8C",x"2D",x"89",x"3B",x"A2",x"B6",x"56",x"09",x"CB",x"E6",x"08",x"D6",x"82",x"B5",x"94",x"B9",x"29",x"38",x"0F",x"09",x"6F",x"E3",x"E6",x"68",x"3C",x"D5",x"AD",x"AB",x"9B",x"82",x"8E",x"30",x"B3",x"AE",x"6E",x"89",x"3A",x"D2",x"4D",x"D2",x"89",x"C9",x"BB",x"32",x"65",x"6B",x"CB",x"56",x"DC",x"5D",x"2C",x"DC",x"12",x"DD",x"F0",x"F1",x"00",x"FF",
		x"60",x"A2",x"2B",x"98",x"3A",x"2B",x"62",x"87",x"B6",x"18",x"52",x"EE",x"5C",x"DC",x"8A",x"92",x"49",x"39",x"75",x"53",x"CA",x"42",x"E0",x"54",x"8D",x"8D",x"2E",x"B3",x"5D",x"24",x"A2",x"1A",x"0B",x"C0",x"15",x"C9",x"16",x"C5",x"22",x"EE",x"31",x"B1",x"47",x"98",x"B2",x"BA",x"FB",x"4E",x"1E",x"61",x"C8",x"C9",x"53",x"5D",x"78",x"24",x"21",x"25",x"F5",x"54",x"E5",x"92",x"07",x"1B",x"11",x"DC",x"53",x"42",x"96",x"7C",x"98",x"92",x"D7",x"0D",x"49",x"74",x"E1",x"E6",x"99",x"34",x"C4",x"39",x"B8",x"A9",x"45",x"93",x"14",x"66",x"6F",x"E1",x"91",x"8D",x"43",x"18",x"43",x"6A",x"54",x"D7",x"0E",x"71",x"F4",x"69",x"11",x"9D",x"26",x"24",x"45",x"BB",x"25",x"67",x"5C",x"02",x"F8",x"E9",x"51",x"FA",x"58",x"B2",x"31",x"A6",x"CE",x"E8",x"8B",x"8D",x"71",x"F6",x"26",x"A3",x"2B",x"3A",x"3B",x"59",x"E7",x"8E",x"36",x"CB",x"A9",x"10",x"7D",x"3C",x"9A",x"2C",x"AF",x"4C",x"6C",x"D5",x"A8",x"A2",x"DE",x"54",x"B2",x"45",x"AD",x"08",x"76",x"42",x"39",x"1A",x"97",x"3C",x"84",x"48",x"D2",x"72",x"5C",x"B2",x"94",x"3C",x"90",x"D3",x"49",x"C9",x"B2",x"F1",x"14",x"B4",x"2A",x"29",x"4F",x"B2",x"C2",x"58",x"26",x"A7",x"32",x"89",x"71",x"61",x"99",x"15",x"AA",x"60",x"DA",x"94",x"25",x"49",x"29",x"BC",x"C9",x"2C",x"96",x"C6",x"A3",x"CA",x"A2",x"AB",x"44",x"56",x"8F",x"AA",x"E8",x"CA",x"E0",x"68",x"3C",x"AA",x"6A",x"23",x"4C",x"A3",x"D5",x"A8",x"6A",x"30",x"D3",x"C8",x"D5",x"A3",x"AA",x"4E",x"44",x"B3",x"17",x"A7",x"A6",x"46",x"16",x"8A",x"AE",x"84",x"2A",x"D0",x"3A",x"5D",x"34",x"B6",x"00",x"7A",x"90",x"14",x"40",x"F7",x"E6",x"0C",x"C8",x"41",x"3C",x"55",x"25",x"A4",x"A9",x"59",x"9D",x"12",x"FB",x"28",x"91",x"15",x"69",x"5B",x"18",x"13",x"55",x"44",x"2E",x"1A",x"71",x"4E",x"A2",x"11",x"39",x"6B",x"C4",x"39",x"B0",x"46",x"F6",x"E2",x"91",x"D4",x"C0",x"62",x"D9",x"AB",x"47",x"DE",x"BC",x"08",x"67",x"2D",x"69",x"75",x"0B",x"A2",x"A8",x"B1",x"44",x"00",x"23",x"0B",x"97",x"A5",x"7A",x"51",x"8B",x"4A",x"9A",x"86",x"14",x"D8",x"3C",x"A3",x"51",x"19",x"72",x"41",x"8B",x"C8",x"A6",x"65",x"CE",x"99",x"D5",x"D2",x"D3",x"A5",x"25",x"47",x"55",x"09",x"6F",x"96",x"B6",x"14",x"C4",x"A4",x"2A",x"59",x"58",x"53",x"65",x"B3",x"CC",x"A4",x"66",x"49",x"5E",x"CD",x"23",x"DB",x"B8",x"23",x"77",x"56",x"77",x"4B",x"43",x"56",x"9B",x"A1",x"DA",x"22",x"C6",x"03",x"FF",
		x"60",x"02",x"A8",x"D9",x"54",x"01",x"35",x"87",x"29",x"A0",x"D5",x"8C",x"D4",x"C5",x"24",x"6E",x"6E",x"89",x"4B",x"E3",x"07",x"B5",x"46",x"B6",x"6A",x"55",x"AC",x"DA",x"EA",x"BE",x"64",x"D4",x"C9",x"55",x"85",x"FA",x"DC",x"51",x"67",x"D7",x"15",x"9C",x"73",x"47",x"9D",x"7C",x"A7",x"4B",x"CD",x"1D",x"75",x"76",x"9D",x"2E",x"35",x"67",x"34",x"39",x"56",x"98",x"75",x"9D",x"D5",x"E6",x"90",x"61",x"5E",x"8D",x"57",x"57",x"7D",x"B8",x"47",x"CE",x"5E",x"5D",x"75",x"6E",x"9E",x"39",x"67",x"F5",x"D5",x"B9",x"78",x"55",x"95",x"D5",x"57",x"6D",x"1C",x"55",x"65",x"57",x"5F",x"8D",x"89",x"7B",x"44",x"6B",x"73",x"8E",x"E5",x"E6",x"5D",x"7B",x"74",x"D5",x"87",x"BB",x"E7",x"EC",x"D1",x"55",x"E7",x"E6",x"99",x"73",x"5A",x"5F",x"9D",x"89",x"57",x"CF",x"69",x"69",x"B1",x"2A",x"9E",x"55",x"65",x"44",x"39",x"B0",x"59",x"4D",x"9C",x"11",x"64",x"27",x"E6",x"B1",x"B1",x"4B",x"18",x"B5",x"96",x"D7",x"58",x"2E",x"F1",x"D6",x"69",x"6A",x"12",x"DB",x"00",x"93",x"BA",x"2A",x"60",x"20",x"97",x"12",x"75",x"9E",x"22",x"9E",x"AB",x"5A",x"D0",x"AC",x"B3",x"47",x"B4",x"0E",x"61",x"73",x"64",x"15",x"99",x"C4",x"B5",x"89",x"84",x"97",x"59",x"DC",x"30",x"46",x"54",x"E9",x"6E",x"71",x"D3",x"E0",x"65",x"BB",x"69",x"2D",x"69",x"63",x"88",x"E1",x"9A",x"5B",x"76",x"8C",x"59",x"B7",x"AB",x"D6",x"95",x"31",x"16",x"5D",x"6E",x"9A",x"77",x"C6",x"94",x"65",x"45",x"88",x"5F",x"09",x"4B",x"34",x"15",x"4E",x"7E",x"55",x"ED",x"5E",x"55",x"9A",x"78",x"9D",x"34",x"05",x"9F",x"43",x"3C",x"51",x"DB",x"E4",x"D2",x"98",x"66",x"86",x"6B",x"B3",x"F7",x"6B",x"16",x"15",x"B4",x"CD",x"DE",x"5C",x"BA",x"7A",x"E5",x"B4",x"58",x"B7",x"A1",x"9C",x"71",x"CD",x"EA",x"E4",x"98",x"4B",x"38",x"31",x"8B",x"B1",x"59",x"42",x"15",x"C5",x"CC",x"CE",x"55",x"19",x"45",x"95",x"36",x"15",x"EB",x"25",x"DC",x"B3",x"DB",x"92",x"43",x"14",x"C5",x"C4",x"6A",x"4B",x"CA",x"91",x"D4",x"1D",x"B9",x"AD",x"A9",x"46",x"D2",x"B6",x"ED",x"B1",x"A6",x"14",x"4D",x"DD",x"71",x"DA",x"96",x"52",x"0C",x"E7",x"C4",x"69",x"7B",x"CA",x"D9",x"54",x"13",x"A5",x"6D",x"B1",x"47",x"6A",x"4E",x"95",x"B2",x"C5",x"96",x"A9",x"D9",x"51",x"D3",x"16",x"96",x"87",x"F6",x"C4",x"6D",x"7B",x"B6",x"D9",x"29",x"3E",x"A5",x"6D",x"59",x"65",x"B7",x"F0",x"D3",x"B0",x"C6",x"DC",x"69",x"5A",x"63",x"CD",x"E1",x"CB",x"98",x"67",x"55",x"31",x"7B",x"E8",x"E9",x"EA",x"1D",x"C6",x"ED",x"D1",x"66",x"3B",x"C6",x"64",x"77",x"44",x"3B",x"1D",x"CC",x"73",x"D4",x"1E",x"5D",x"97",x"A1",x"4D",x"7D",x"FF",
		x"60",x"6C",x"D2",x"6A",x"D2",x"45",x"EC",x"AA",x"8E",x"B7",x"56",x"56",x"4F",x"52",x"1A",x"E7",x"26",x"93",x"B1",x"49",x"AB",x"9C",x"3B",x"37",x"E5",x"D5",x"A3",x"0C",x"EA",x"43",x"4D",x"3A",x"B7",x"32",x"C4",x"D5",x"54",x"EE",x"55",x"4A",x"DF",x"43",x"4B",x"64",x"55",x"A9",x"C2",x"54",x"2D",x"95",x"D5",x"A5",x"0E",x"83",x"B2",x"58",x"DB",x"A4",x"36",x"6E",x"8A",x"10",x"5E",x"93",x"FA",x"B2",x"C9",x"CD",x"78",x"73",x"1B",x"9B",x"0B",x"83",x"CC",x"C6",x"63",x"EA",x"C6",x"8D",x"3C",x"2B",x"B5",x"A9",x"79",x"57",x"CA",x"2C",x"D5",x"A6",x"92",x"45",x"B5",x"BC",x"52",x"9B",x"4B",x"11",x"F1",x"F2",x"2E",x"E5",x"C8",x"43",x"25",x"9C",x"DB",x"A6",x"2D",x"0F",x"B6",x"52",x"59",x"13",x"8E",x"34",x"D0",x"4B",x"6D",x"4B",x"58",x"F3",x"34",x"F5",x"A4",x"76",x"61",x"4F",x"39",x"95",x"CB",x"92",x"87",x"33",x"0D",x"11",x"2B",x"4D",x"67",x"F6",x"D4",x"D8",x"C2",x"3D",x"2D",x"DA",x"43",x"85",x"4E",x"F7",x"5A",x"0F",x"FF",
		x"60",x"66",x"4A",x"59",x"8D",x"25",x"1A",x"AB",x"31",x"65",x"75",x"D6",x"6C",x"92",x"86",x"98",x"34",x"D8",x"AB",x"4E",x"A9",x"53",x"F2",x"C2",x"E8",x"25",x"A3",x"2F",x"D6",x"46",x"34",x"D7",x"8C",x"AE",x"58",x"1F",x"95",x"58",x"3B",x"9A",x"A2",x"63",x"8C",x"72",x"C9",x"A8",x"93",x"AD",x"51",x"EA",x"25",x"A3",x"CE",x"AA",x"26",x"20",x"E7",x"8C",x"26",x"C9",x"6A",x"C7",x"BA",x"33",x"EA",x"CC",x"27",x"1C",x"7D",x"09",x"30",x"20",x"45",x"D2",x"D2",x"16",x"13",x"A3",x"92",x"4B",x"5A",x"9D",x"6D",x"B4",x"59",x"39",x"6B",x"79",x"F2",x"11",x"12",x"29",x"AF",x"94",x"A9",x"89",x"58",x"98",x"B6",x"52",x"C6",x"E8",x"E4",x"19",x"EA",x"4B",x"1E",x"12",x"F3",x"86",x"A5",x"2D",x"99",x"0F",x"EC",x"9B",x"D1",x"6A",x"64",x"D9",x"88",x"46",x"57",x"A6",x"96",x"25",x"A9",x"1E",x"5B",x"0D",x"46",x"5A",x"AD",x"88",x"74",x"4F",x"1C",x"49",x"37",x"C6",x"14",x"39",x"7B",x"24",x"C3",x"1A",x"93",x"C7",x"94",x"11",x"36",x"2B",x"24",x"5D",x"53",x"46",x"50",x"15",x"73",x"74",x"D7",x"6D",x"41",x"33",x"24",x"5E",x"5D",x"2F",x"85",x"C5",x"A0",x"56",x"E7",x"D4",x"10",x"65",x"41",x"D9",x"95",x"A1",x"42",x"54",x"2D",x"B3",x"56",x"16",x"4A",x"49",x"B3",x"CA",x"1C",x"55",x"39",x"C4",x"5D",x"2B",x"73",x"44",x"19",x"17",x"56",x"C7",x"64",x"95",x"75",x"4D",x"50",x"15",x"B3",x"55",x"CD",x"53",x"41",x"D1",x"A4",x"51",x"55",x"8F",x"87",x"0F",x"FF",
		x"60",x"6A",x"E5",x"76",x"D3",x"44",x"9C",x"A8",x"95",x"97",x"76",x"13",x"71",x"1A",x"16",x"15",x"2B",x"4C",x"29",x"75",x"59",x"5C",x"71",x"D5",x"F0",x"CD",x"6D",x"4D",x"41",x"C2",x"C2",x"1E",x"8D",x"A5",x"06",x"53",x"0E",x"5F",x"3B",x"E6",x"66",x"4C",x"29",x"F2",x"C9",x"98",x"BB",x"35",x"67",x"D6",x"27",x"65",x"C9",x"5A",x"4D",x"E5",x"2A",x"B7",x"A5",x"D1",x"94",x"50",x"9F",x"A4",x"80",x"C9",x"CB",x"47",x"5F",x"8D",x"9B",x"70",x"2C",x"19",x"6D",x"F6",x"6A",x"EC",x"D5",x"64",x"D4",x"39",x"29",x"5B",x"44",x"E7",x"51",x"E6",x"A6",x"14",x"A1",x"BD",x"5A",x"96",x"2B",x"71",x"85",x"F6",x"6E",x"49",x"EE",x"44",x"95",x"DA",x"AB",x"C4",x"65",x"A3",x"A4",x"DA",x"A6",x"12",x"95",x"86",x"6A",x"19",x"99",x"53",x"94",x"83",x"8A",x"79",x"B4",x"4A",x"61",x"2E",x"4A",x"1E",x"96",x"39",x"C4",x"25",x"A9",x"72",x"84",x"DB",x"14",x"65",x"A9",x"66",x"59",x"B6",x"5D",x"9C",x"2B",x"53",x"A4",x"A5",x"21",x"51",x"69",x"C2",x"9C",x"69",x"EF",x"01",x"FF",
		x"60",x"25",x"CF",x"D6",x"22",x"BA",x"2A",x"8F",x"AC",x"78",x"D3",x"E8",x"9C",x"3C",x"92",x"12",x"CD",x"2C",x"BA",x"F1",x"88",x"B3",x"6E",x"73",x"AB",x"D9",x"23",x"89",x"FA",x"5C",x"B4",x"A7",x"8C",x"2C",x"8A",x"4B",x"A3",x"9E",x"32",x"F2",x"8C",x"AF",x"83",x"AC",x"6E",x"CB",x"13",x"B9",x"2E",x"F4",x"BA",x"A5",x"08",x"7C",x"3B",x"39",x"EC",x"85",x"C4",x"7B",x"F3",x"9A",x"30",x"5D",x"E2",x"1C",x"5C",x"3D",x"BB",x"4E",x"89",x"93",x"19",x"B3",x"A8",x"39",x"25",x"C9",x"62",x"32",x"34",x"93",x"A5",x"3C",x"F1",x"C9",x"D2",x"88",x"9A",x"DA",x"42",x"3A",x"CB",x"22",x"8A",x"2B",x"12",x"EB",x"6C",x"4B",x"A9",x"04",x"D0",x"7E",x"1C",x"01",x"5E",x"79",x"20",x"A0",x"CB",x"30",x"02",x"24",x"17",x"86",x"80",x"A4",x"23",x"10",x"E0",x"5D",x"26",x"02",x"AC",x"F0",x"78",x"FF",
		x"60",x"2A",x"10",x"79",x"4C",x"C5",x"92",x"04",x"D7",x"4D",x"65",x"AB",x"58",x"59",x"9C",x"D8",x"5C",x"B4",x"A3",x"41",x"71",x"7D",x"71",x"CF",x"EA",x"C9",x"CD",x"0D",x"D5",x"B5",x"AA",x"AD",x"36",x"2F",x"A4",x"A1",x"AC",x"09",x"D7",x"BC",x"E0",x"8F",x"3C",x"B7",x"6A",x"F3",x"82",x"78",x"17",x"A9",x"A9",x"25",x"B0",x"E6",x"43",x"34",x"EB",x"A6",x"34",x"A2",x"2F",x"51",x"6F",x"1C",x"BA",x"D8",x"82",x"9D",x"33",x"B1",x"EB",x"43",x"36",x"8F",x"EC",x"99",x"AA",x"F7",x"D5",x"AD",x"AA",x"E3",x"2A",x"A0",x"74",x"93",x"56",x"04",x"9F",x"D2",x"5E",x"76",x"46",x"9B",x"74",x"B9",x"46",x"2C",x"1A",x"7D",x"96",x"5D",x"A2",x"BE",x"69",x"0C",x"59",x"74",x"8B",x"DA",x"EA",x"31",x"16",x"5E",x"2D",x"66",x"AB",x"DA",x"9C",x"EC",x"06",x"BA",x"2F",x"6E",x"6B",x"A3",x"51",x"E2",x"DC",x"24",x"AD",x"C5",x"A8",x"0B",x"85",x"DD",x"B0",x"55",x"A1",x"66",x"6C",x"75",x"C3",x"96",x"65",x"BA",x"69",x"D4",x"09",x"5B",x"E1",x"91",x"AE",x"D6",x"38",x"EC",x"45",x"64",x"99",x"58",x"13",x"33",x"16",x"9E",x"2D",x"6A",x"B3",x"CC",x"9C",x"75",x"A7",x"A8",x"D5",x"11",x"7B",x"A5",x"51",x"A2",x"92",x"F8",x"01",x"FF",
		x"60",x"6D",x"6C",x"5E",x"93",x"3B",x"97",x"B4",x"39",x"7B",x"29",x"DD",x"AE",x"3D",x"A6",x"E2",x"35",x"B9",x"73",x"F6",x"18",x"B3",x"F5",x"A6",x"AE",x"D9",x"A3",x"CF",x"3A",x"47",x"B9",x"E6",x"8C",x"3A",x"CA",x"6B",x"15",x"9F",x"55",x"6A",x"E7",x"BE",x"14",x"6B",x"6A",x"09",x"54",x"7A",x"63",x"E9",x"A8",x"C9",x"37",x"E5",x"54",x"29",x"94",x"A6",x"26",x"1B",x"37",x"F7",x"B6",x"5D",x"CA",x"66",x"3C",x"5D",x"33",x"49",x"19",x"AB",x"F2",x"0A",x"CD",x"26",x"A5",x"2B",x"32",x"2B",x"34",x"E2",x"85",x"38",x"A8",x"4D",x"F7",x"B0",x"EB",x"62",x"6F",x"36",x"93",x"CD",x"9E",x"0B",x"BC",x"DE",x"2C",x"73",x"3A",x"CE",x"CF",x"3C",x"22",x"3D",x"62",x"09",x"A0",x"F8",x"54",x"02",x"F8",x"14",x"4E",x"00",x"E7",x"5D",x"11",x"E0",x"4D",x"E8",x"03",x"FF",
		x"60",x"AA",x"0E",x"5C",x"2A",x"CD",x"63",x"9B",x"39",x"28",x"29",x"B3",x"B2",x"9C",x"C6",x"A6",x"D0",x"32",x"AD",x"72",x"1B",x"67",x"14",x"23",x"F3",x"C7",x"6D",x"5A",x"49",x"1D",x"C5",x"9E",x"8C",x"79",x"27",x"33",x"64",x"5D",x"33",x"E6",x"15",x"C3",x"81",x"74",x"CD",x"98",x"57",x"74",x"43",x"92",x"37",x"66",x"AB",x"9C",x"45",x"2D",x"67",x"21",x"00",x"84",x"6C",x"05",x"04",x"61",x"61",x"80",x"4A",x"D5",x"0C",x"D0",x"AD",x"29",x"03",x"0A",x"65",x"67",x"40",x"A6",x"EC",x"04",x"48",x"5C",x"CC",x"E4",x"C5",x"B8",x"B9",x"99",x"93",x"90",x"FB",x"A4",x"61",x"9C",x"AB",x"5B",x"16",x"7C",x"58",x"B0",x"77",x"29",x"51",x"F0",x"E1",x"CE",x"D6",x"A5",x"04",x"CE",x"87",x"07",x"7B",x"E6",x"12",x"38",x"5F",x"12",x"14",x"9D",x"4A",x"EC",x"D5",x"58",x"AA",x"64",x"2A",x"99",x"B7",x"A5",x"89",x"DA",x"39",x"15",x"4E",x"B5",x"15",x"4B",x"A7",x"54",x"5B",x"9B",x"56",x"A4",x"9D",x"53",x"E3",x"65",x"6B",x"B1",x"B6",x"49",x"43",x"E4",x"29",x"C3",x"92",x"26",x"4C",x"D1",x"8B",x"14",x"7B",x"6A",x"33",x"7B",x"57",x"9A",x"E4",x"A9",x"C3",x"56",x"8D",x"9B",x"45",x"48",x"31",x"79",x"34",x"AA",x"19",x"29",x"D5",x"94",x"41",x"79",x"A4",x"85",x"15",x"55",x"07",x"63",x"56",x"E1",x"B6",x"45",x"EB",x"45",x"59",x"9A",x"B9",x"01",x"00",x"00",x"37",x"55",x"EF",x"6E",x"6C",x"B1",x"5B",x"9B",x"2B",x"B9",x"77",x"CE",x"1D",x"6D",x"49",x"1A",x"52",x"39",x"67",x"54",x"B5",x"78",x"72",x"C6",x"DC",x"91",x"97",x"64",x"A1",x"55",x"4B",x"46",x"5A",x"B2",x"A5",x"56",x"D5",x"19",x"51",x"C9",x"9A",x"3A",x"5D",x"67",x"84",x"29",x"49",x"C6",x"54",x"9C",x"11",x"E6",x"24",x"21",x"D7",x"B6",x"53",x"92",x"BD",x"BA",x"7A",x"35",x"86",x"56",x"D5",x"E4",x"21",x"1E",x"31",x"47",x"5D",x"7C",x"A8",x"5B",x"46",x"1C",x"6D",x"F1",x"21",x"61",x"15",x"69",x"75",x"C5",x"9B",x"8B",x"6D",x"E4",x"31",x"94",x"C4",x"1A",x"DD",x"51",x"DA",x"54",x"22",x"8B",x"76",x"D5",x"4B",x"4B",x"D1",x"14",x"36",x"5B",x"25",x"6D",x"CD",x"B0",x"68",x"F5",x"54",x"73",x"14",x"49",x"16",x"D9",x"71",x"1F",x"FF",
		x"60",x"69",x"4C",x"C9",x"5C",x"35",x"EB",x"B4",x"31",x"25",x"4B",x"8E",x"99",x"DB",x"86",x"1C",x"BD",x"29",x"6B",x"49",x"EB",x"72",x"88",x"C1",x"8A",x"B9",x"AD",x"2D",x"C6",x"97",x"DC",x"E7",x"B6",x"AA",x"48",x"3B",x"36",x"BF",x"DD",x"F2",x"24",x"73",x"85",x"6A",x"55",x"CB",x"33",x"9E",x"4A",x"F4",x"D5",x"A5",x"CC",x"34",x"CB",x"D9",x"32",x"03",x"01",x"62",x"D5",x"64",x"40",x"6C",x"96",x"A5",x"28",x"21",x"9A",x"2A",x"92",x"94",x"3A",x"99",x"68",x"2C",x"B5",x"DB",x"86",x"18",x"DC",x"B8",x"55",x"6B",x"19",x"63",x"0E",x"4A",x"77",x"6D",x"69",x"8A",x"85",x"A5",x"4C",x"B3",x"A6",x"29",x"37",x"4C",x"B3",x"D8",x"D4",x"96",x"52",x"58",x"A5",x"6C",x"F5",x"58",x"9A",x"77",x"C5",x"F0",x"35",x"63",x"9D",x"DA",x"0C",x"3D",x"96",x"B4",x"B5",x"6B",x"13",x"F6",x"5C",x"DC",x"96",x"6E",x"4D",x"C4",x"AA",x"EE",x"98",x"9B",x"77",x"26",x"EB",x"38",x"6D",x"6A",x"52",x"C4",x"62",x"1B",x"B7",x"B1",x"19",x"65",x"F1",x"6D",x"D4",x"86",x"E6",x"94",x"C5",x"27",x"71",x"EA",x"B3",x"66",x"B5",x"ED",x"44",x"A9",x"CF",x"42",x"C2",x"B7",x"62",x"86",x"BE",x"18",x"11",x"ED",x"AE",x"AD",x"E6",x"96",x"CD",x"D0",x"32",x"B1",x"19",x"5B",x"76",x"25",x"CD",x"24",x"66",x"6C",x"46",x"59",x"7C",x"1B",x"99",x"A1",x"39",x"65",x"F1",x"49",x"2C",x"FA",x"AC",x"59",x"6D",x"3B",x"91",x"E8",x"B3",x"90",x"F0",x"AD",x"98",x"0F",x"FF",
		x"60",x"6C",x"D6",x"76",x"2A",x"44",x"EC",x"8A",x"45",x"FA",x"0D",x"17",x"76",x"2A",x"16",x"E5",x"36",x"CC",x"44",x"89",x"5A",x"45",x"1C",x"77",x"16",x"3B",x"6E",x"96",x"B9",x"C3",x"49",x"92",x"94",x"D1",x"E5",x"48",x"56",x"EB",x"3A",x"BA",x"9C",x"2C",x"C4",x"A4",x"EB",x"A8",x"6A",x"0C",x"56",x"B5",x"75",x"A3",x"E8",x"32",x"44",x"CC",x"5E",x"8D",x"B2",x"DA",x"10",x"E1",x"B8",x"5D",x"BA",x"C1",x"4C",x"35",x"6C",x"A1",x"00",x"96",x"28",x"2B",x"63",x"51",x"61",x"6A",x"31",x"6B",x"0C",x"D9",x"AB",x"73",x"C6",x"DC",x"31",x"16",x"A3",x"26",x"6D",x"5D",x"C6",x"58",x"92",x"B2",x"A7",x"B5",x"1B",x"63",x"C9",x"46",x"9E",x"DA",x"6E",x"0C",x"A5",x"19",x"79",x"51",x"97",x"D6",x"97",x"A9",x"EC",x"81",x"7D",x"5A",x"5F",x"86",x"90",x"27",x"F7",x"19",x"5D",x"E9",x"42",x"1E",x"DA",x"75",x"74",x"25",x"1B",x"49",x"44",x"96",x"D0",x"A4",x"40",x"66",x"19",x"A9",x"C3",x"90",x"23",x"73",x"A6",x"B6",x"76",x"43",x"C9",x"CE",x"9A",x"92",x"34",x"0C",x"D9",x"A9",x"72",x"8E",x"D3",x"D0",x"E5",x"28",x"CA",x"5D",x"C9",x"4C",x"57",x"9A",x"90",x"A5",x"67",x"65",x"5D",x"A9",x"4A",x"1A",x"91",x"E5",x"01",x"FF",
		x"60",x"AC",x"52",x"72",x"22",x"CC",x"EC",x"A8",x"5C",x"A6",x"36",x"33",x"B3",x"93",x"22",x"5B",x"DC",x"4C",x"AC",x"F3",x"08",x"42",x"94",x"08",x"8B",x"85",x"23",x"C8",x"5E",x"29",x"BD",x"1A",x"8D",x"A8",x"6A",x"67",x"93",x"5C",x"D4",x"F2",x"CE",x"93",x"9D",x"6D",x"B1",x"00",x"86",x"28",x"69",x"DD",x"10",x"29",x"C6",x"D2",x"68",x"54",x"C5",x"BA",x"88",x"C6",x"9C",x"51",x"57",x"E3",x"2A",x"66",x"6B",x"46",x"57",x"A2",x"B3",x"B8",x"AF",x"19",x"43",x"49",x"2E",x"DC",x"DE",x"75",x"8C",x"39",x"2A",x"6B",x"7B",x"9F",x"31",x"E5",x"A8",x"6C",x"ED",x"79",x"C6",x"94",x"92",x"70",x"54",x"74",x"19",x"73",x"0A",x"CA",x"51",x"D1",x"6E",x"CC",x"39",x"0B",x"47",x"58",x"D7",x"B1",x"E4",x"C2",x"12",x"A1",x"5D",x"C7",x"9A",x"0B",x"8B",x"A7",x"74",x"1D",x"5B",x"49",x"2E",x"54",x"D2",x"B7",x"6D",x"D9",x"A8",x"61",x"47",x"9B",x"B4",x"17",x"A3",x"81",x"51",x"4D",x"DD",x"91",x"32",x"73",x"A4",x"75",x"71",x"47",x"AE",x"2C",x"E1",x"DA",x"D5",x"2D",x"25",x"2B",x"7B",x"48",x"5A",x"B3",x"15",x"E3",x"2C",x"9E",x"C9",x"CC",x"16",x"95",x"8B",x"CF",x"4C",x"12",x"7B",x"54",x"66",x"5E",x"53",x"F9",x"01",x"FF",
		x"60",x"6A",x"E9",x"0C",x"CD",x"A3",x"2A",x"A7",x"B1",x"05",x"32",x"CC",x"5A",x"5C",x"86",x"14",x"28",x"34",x"62",x"71",x"EA",x"42",x"96",x"50",x"8F",x"2D",x"69",x"0A",x"55",x"53",x"D4",x"37",x"A7",x"29",x"34",x"2D",x"56",x"DF",x"9C",x"A6",x"D8",x"A4",x"44",x"63",x"73",x"99",x"52",x"95",x"12",x"B7",x"CD",x"65",x"49",x"59",x"42",x"5A",x"37",x"97",x"36",x"39",x"49",x"CE",x"CC",x"53",x"BA",x"A2",x"A5",x"21",x"B2",x"57",x"99",x"8A",x"E2",x"41",x"ED",x"4E",x"61",x"8A",x"C6",x"1A",x"A5",x"9B",x"B4",x"31",x"E4",x"4E",x"CA",x"9A",x"33",x"FA",x"14",x"BA",x"D9",x"AB",x"E9",x"E8",x"4A",x"88",x"51",x"AB",x"35",x"A3",x"AE",x"3E",x"DD",x"22",x"D7",x"8C",x"BC",x"38",x"51",x"AF",x"A9",x"3C",x"F2",x"A6",x"95",x"A5",x"7A",x"4E",x"2A",x"8B",x"03",x"8F",x"AA",x"28",x"02",x"A8",x"31",x"42",x"00",x"D5",x"65",x"86",x"AE",x"F8",x"2C",x"B7",x"68",x"2A",x"80",x"1A",x"22",x"4D",x"5E",x"BD",x"AA",x"65",x"CF",x"66",x"40",x"D7",x"C6",x"02",x"70",x"D9",x"3B",x"54",x"BA",x"67",x"1A",x"7A",x"92",x"56",x"D9",x"D8",x"91",x"22",x"49",x"5A",x"E9",x"62",x"5B",x"2B",x"75",x"29",x"85",x"6B",x"C1",x"6D",x"BA",x"39",x"95",x"BE",x"B1",x"B7",x"FA",x"EB",x"54",x"C6",x"8A",x"D1",x"16",x"1B",x"53",x"95",x"0A",x"A6",x"7B",x"36",x"4C",x"75",x"E7",x"1C",x"D9",x"E6",x"88",x"01",x"93",x"68",x"30",x"A0",x"E3",x"34",x"06",x"74",x"D0",x"69",x"8A",x"8A",x"D7",x"82",x"A3",x"A9",x"2A",x"2B",x"59",x"B2",x"CC",x"64",x"AA",x"6C",x"6A",x"C8",x"24",x"92",x"32",x"A0",x"92",x"60",x"02",x"4C",x"95",x"46",x"80",x"C9",x"53",x"CC",x"56",x"B8",x"71",x"54",x"57",x"4E",x"7D",x"56",x"22",x"51",x"3D",x"BA",x"74",x"59",x"98",x"7A",x"E5",x"C4",x"D4",x"17",x"A1",x"52",x"D2",x"0B",x"C3",x"34",x"A5",x"89",x"B8",x"AC",x"62",x"40",x"E4",x"64",x"04",x"F0",x"56",x"14",x"01",x"3E",x"A3",x"99",x"2E",x"3B",x"13",x"33",x"8D",x"6A",x"AA",x"60",x"DC",x"22",x"CC",x"AA",x"2B",x"4D",x"72",x"73",x"4F",x"79",x"25",x"F1",x"95",x"DA",x"B4",x"1A",x"B7",x"38",x"54",x"2B",x"89",x"2A",x"D3",x"E2",x"58",x"25",x"A5",x"3B",x"EA",x"88",x"52",x"92",x"E4",x"8B",x"2A",x"29",x"8C",x"9A",x"87",x"D3",x"65",x"95",x"20",x"1B",x"4E",x"F3",x"96",x"34",x"C2",x"6A",x"C5",x"BC",x"26",x"CC",x"08",x"9B",x"62",x"9B",x"8A",x"B0",x"25",x"4C",x"46",x"2A",x"25",x"AD",x"94",x"30",x"19",x"19",x"09",x"57",x"9C",x"82",x"68",x"A5",x"A4",x"C3",x"56",x"B1",x"4B",x"E0",x"D2",x"EE",x"DA",x"2A",x"4C",x"41",x"52",x"A3",x"4D",x"A5",x"B0",x"78",x"75",x"F3",x"50",x"D6",x"AA",x"DC",x"C3",x"C3",x"B2",x"4A",x"CB",x"D2",x"74",x"77",x"AF",x"AA",x"2D",x"4F",x"53",x"4B",x"AA",x"A3",x"B6",x"32",x"F6",x"08",x"8B",x"AA",x"32",x"EA",x"98",x"AA",x"CC",x"72",x"D1",x"E8",x"42",x"EC",x"70",x"8D",x"59",x"6D",x"0C",x"A1",x"33",x"28",x"16",x"B7",x"D9",x"A7",x"28",x"95",x"4A",x"DC",x"F6",x"58",x"5D",x"C3",x"C2",x"32",x"03",x"C2",x"A0",x"72",x"65",x"EA",x"1E",x"E6",x"55",x"C5",x"D5",x"31",x"55",x"B9",x"E6",x"22",x"D3",x"86",x"58",x"69",x"9A",x"8B",x"D4",x"10",x"7C",x"55",x"51",x"2C",x"66",x"40",x"17",x"E1",x"04",x"88",x"B4",x"93",x"00",x"89",x"87",x"22",x"A0",x"38",x"C7",x"07",x"FF",
		x"60",x"69",x"8C",x"36",x"16",x"C3",x"17",x"A7",x"3E",x"9A",x"38",x"74",x"9F",x"5D",x"BA",x"A4",x"FC",x"44",x"AD",x"75",x"69",x"8A",x"94",x"73",x"95",x"D6",x"AD",x"A9",x"52",x"DB",x"54",x"B7",x"8C",x"BA",x"C8",x"70",x"8E",x"5C",x"D5",x"EA",x"26",x"55",x"29",x"62",x"F5",x"28",x"BB",x"36",x"A1",x"C8",x"46",x"2D",x"AF",x"C1",x"48",x"2A",x"33",x"B7",x"2C",x"06",x"A3",x"8E",x"4A",x"D3",x"B2",x"94",x"D5",x"4A",x"AD",x"4B",x"CB",x"62",x"76",x"F3",x"B0",x"6C",x"C0",x"00",x"19",x"22",x"04",x"10",x"A5",x"7B",x"CA",x"73",x"50",x"4F",x"B3",x"88",x"29",x"CB",x"DE",x"2D",x"C4",x"CB",x"94",x"28",x"75",x"4B",x"F5",x"B6",x"DB",x"C2",x"D8",x"C3",x"32",x"AA",x"6C",x"8B",x"52",x"69",x"F1",x"8C",x"29",x"2D",x"8A",x"AD",x"24",x"32",x"26",x"B7",x"28",x"8C",x"D4",x"CC",x"98",x"DC",x"E2",x"D0",x"3D",x"52",x"62",x"51",x"8B",x"43",x"D3",x"68",x"91",x"D5",x"25",x"09",x"8D",x"A3",x"45",x"DA",x"94",x"34",x"4E",x"F2",x"12",x"6B",x"5A",x"D2",x"34",x"C9",x"5B",x"6C",x"75",x"CB",x"62",x"A3",x"28",x"F5",x"26",x"2D",x"8B",x"8D",x"A2",x"A4",x"6A",x"8F",x"2C",x"F9",x"A4",x"B4",x"68",x"D2",x"F2",x"E4",x"CD",x"D4",x"3A",x"6A",x"A9",x"2B",x"AB",x"30",x"D7",x"D8",x"02",x"C8",x"BA",x"3D",x"34",x"A9",x"B8",x"5A",x"A8",x"53",x"97",x"FB",x"C2",x"51",x"A1",x"49",x"4A",x"E6",x"A2",x"87",x"85",x"B5",x"19",x"69",x"D2",x"16",x"29",x"B6",x"A6",x"A5",x"49",x"67",x"06",x"DB",x"22",x"94",x"47",x"1A",x"AE",x"A6",x"AD",x"4B",x"DA",x"BC",x"9B",x"B8",x"64",x"1A",x"49",x"33",x"CE",x"EC",x"B9",x"AA",x"25",x"CD",x"3A",x"51",x"D4",x"A2",x"91",x"34",x"E7",x"CC",x"96",x"B3",x"47",x"DA",x"98",x"9B",x"AA",x"B7",x"1E",x"49",x"C5",x"A3",x"98",x"D9",x"68",x"C4",x"95",x"AC",x"B1",x"FB",x"A2",x"11",x"25",x"BD",x"6E",x"92",x"B3",x"46",x"18",x"DD",x"B9",x"69",x"2C",x"1E",x"61",x"88",x"EB",x"AE",x"31",x"A7",x"85",x"A1",x"4C",x"B8",x"D4",x"9C",x"16",x"87",x"DA",x"EE",x"DA",x"93",x"5B",x"1A",x"46",x"69",x"D8",x"54",x"69",x"79",x"18",x"69",x"E1",x"53",x"BB",x"15",x"B1",x"94",x"BB",x"D7",x"6C",x"02",x"B8",x"E1",x"46",x"80",x"68",x"37",x"18",x"10",x"ED",x"05",x"01",x"A2",x"BB",x"60",x"40",x"52",x"EF",x"04",x"48",x"E6",x"1C",x"08",x"10",x"B5",x"1B",x"02",x"2A",x"31",x"79",x"FF",
		x"60",x"61",x"CA",x"9A",x"CD",x"7A",x"2A",x"95",x"BA",x"48",x"CC",x"CC",x"AC",x"D4",x"CA",x"C4",x"25",x"CA",x"AB",x"56",x"AA",x"AA",x"70",x"0E",x"CD",x"49",x"0C",x"E8",x"DC",x"38",x"A5",x"85",x"85",x"84",x"D6",x"A4",x"16",x"F9",x"A8",x"5E",x"B9",x"56",x"47",x"12",x"82",x"86",x"FA",x"94",x"75",x"65",x"34",x"EE",x"2A",x"1E",x"C7",x"54",x"91",x"4B",x"57",x"7A",x"2D",x"54",x"14",x"6D",x"62",x"52",x"95",x"5B",x"EC",x"BB",x"4B",x"66",x"95",x"6D",x"69",x"9C",x"E6",x"5A",x"63",x"A7",x"A5",x"B1",x"65",x"68",x"4C",x"D4",x"96",x"C4",x"1A",x"C9",x"B1",x"51",x"5A",x"14",x"AA",x"25",x"D5",x"86",x"29",x"61",x"88",x"96",x"2C",x"BD",x"38",x"44",x"A1",x"70",x"A0",x"77",x"6A",x"95",x"C6",x"61",x"A1",x"35",x"56",x"54",x"1A",x"5B",x"B8",x"F9",x"C6",x"A1",x"A9",x"00",x"8A",x"89",x"6C",x"51",x"B5",x"A9",x"1E",x"5E",x"25",x"F9",x"DE",x"98",x"BB",x"7B",x"D5",x"E2",x"27",x"47",x"29",x"D5",x"55",x"59",x"6E",x"59",x"78",x"46",x"5A",x"44",x"55",x"93",x"A6",x"E2",x"A1",x"B8",x"46",x"23",x"CA",x"5E",x"D4",x"AA",x"A7",x"8E",x"28",x"66",x"CE",x"CE",x"B4",x"32",x"E2",x"58",x"5D",x"32",x"2B",x"6C",x"8B",x"63",x"0F",x"AE",x"8E",x"A8",x"2D",x"8E",x"4B",x"B5",x"33",x"A3",x"B5",x"24",x"8E",x"E4",x"EA",x"B0",x"DA",x"B2",x"D8",x"43",x"A3",x"2A",x"CC",x"28",x"63",x"0F",x"8D",x"AA",x"B0",x"A3",x"89",x"8B",x"23",x"33",x"EC",x"8C",x"3E",x"76",x"4B",x"ED",x"B6",x"3B",x"86",x"34",x"D5",x"BD",x"DB",x"EE",x"98",x"52",x"B5",x"92",x"1A",x"3B",x"6D",x"89",x"5D",x"33",x"33",x"A3",x"94",x"35",x"16",x"2D",x"EF",x"96",x"9B",x"F6",x"50",x"B5",x"2A",x"CB",x"6E",x"38",x"62",x"B1",x"CC",x"CC",x"78",x"E1",x"48",x"D9",x"22",x"32",x"E2",x"B9",x"BD",x"44",x"75",x"CB",x"8C",x"6B",x"F6",x"1A",x"38",x"A4",x"4B",x"8A",x"D9",x"5B",x"64",x"E3",x"9E",x"3A",x"0F",x"FF",
		x"60",x"26",x"B2",x"7A",x"4C",x"A4",x"1B",x"87",x"20",x"13",x"CD",x"16",x"EB",x"3A",x"BC",x"E2",x"DD",x"85",x"37",x"C9",x"F2",x"B3",x"33",x"D7",x"9C",x"DA",x"2B",x"2A",x"CE",x"42",x"72",x"EA",x"8C",x"B8",x"86",x"30",x"96",x"9E",x"AA",x"AA",x"28",x"4D",x"25",x"3A",x"0A",x"08",x"A0",x"EA",x"34",x"05",x"64",x"13",x"E6",x"A2",x"E2",x"DC",x"D5",x"A6",x"89",x"8B",x"9B",x"0B",x"17",x"CE",x"39",x"0C",x"E8",x"D0",x"85",x"01",x"9D",x"BB",x"30",x"60",x"30",x"E7",x"94",x"36",x"63",x"2C",x"9A",x"B5",x"5B",x"DC",x"AD",x"31",x"6A",x"DD",x"69",x"E9",x"52",x"2C",x"A2",x"75",x"A7",x"E4",x"4B",x"B3",x"90",x"CE",x"E3",x"92",x"6F",x"4D",x"C2",x"3A",x"8B",x"53",x"B1",x"15",x"8A",x"DA",x"2C",x"49",x"C5",x"B6",x"24",x"AC",x"BD",x"BA",x"E5",x"C3",x"A9",x"80",x"55",x"EB",x"96",x"17",x"CF",x"62",x"15",x"5D",x"4A",x"E1",x"AD",x"46",x"7A",x"74",x"49",x"65",x"50",x"95",x"62",x"9E",x"37",x"94",x"49",x"75",x"A2",x"A9",x"1B",x"54",x"55",x"EE",x"49",x"62",x"4E",x"4B",x"D3",x"72",x"85",x"06",x"DB",x"19",x"55",x"CB",x"22",x"92",x"DE",x"65",x"34",x"35",x"AA",x"69",x"C4",x"9A",x"D1",x"55",x"A7",x"AE",x"1E",x"4F",x"C4",x"D0",x"BC",x"BB",x"0A",x"2E",x"19",x"5D",x"35",x"1A",x"1A",x"7E",x"7B",x"74",x"C5",x"79",x"AA",x"77",x"EB",x"D1",x"16",x"1B",x"19",x"52",x"4D",x"46",x"5B",x"5C",x"66",x"48",x"2D",x"1D",x"5D",x"B6",x"99",x"29",x"35",x"67",x"74",x"C9",x"67",x"B8",x"F5",x"94",x"36",x"64",x"23",x"C3",x"51",x"AD",x"C6",x"50",x"9C",x"16",x"5B",x"35",x"1E",x"7D",x"B1",x"1E",x"AA",x"D9",x"64",x"0C",x"D9",x"86",x"9B",x"66",x"93",x"D6",x"26",x"1B",x"EE",x"5A",x"B5",x"4B",x"97",x"5D",x"7A",x"5A",x"56",x"0D",x"5D",x"B1",x"D2",x"6A",x"D5",x"C4",x"F5",x"C9",x"A8",x"87",x"7B",x"98",x"D4",x"57",x"6B",x"69",x"9A",x"CD",x"D3",x"50",x"95",x"87",x"6B",x"B6",x"63",x"40",x"55",x"E6",x"AD",x"9F",x"5E",x"15",x"2D",x"E7",x"8C",x"6E",x"06",x"57",x"94",x"5C",x"33",x"DA",x"19",x"C2",x"90",x"63",x"CD",x"68",x"47",x"2C",x"43",x"8E",x"AE",x"A3",x"EB",x"21",x"84",x"2C",x"DB",x"8D",x"A1",x"A5",x"10",x"0A",x"5F",x"37",x"C6",x"9A",x"5D",x"B8",x"6C",x"CB",x"98",x"6A",x"71",x"95",x"B4",x"AE",x"63",x"AA",x"D9",x"54",x"CA",x"BA",x"8D",x"B9",x"E4",x"50",x"49",x"4F",x"37",x"96",x"92",x"C3",x"24",x"3C",x"DB",x"58",x"4B",x"75",x"93",x"D0",x"EE",x"6D",x"2D",x"CB",x"DD",x"9C",x"9B",x"A6",x"BD",x"14",x"33",x"4D",x"ED",x"62",x"F6",x"DC",x"D1",x"A3",x"BC",x"A6",x"3A",x"62",x"E4",x"C8",x"F6",x"86",x"EA",x"8A",x"89",x"23",x"CB",x"1B",x"92",x"27",x"16",x"8A",x"18",x"6F",x"F8",x"00",x"FF",
		x"60",x"C5",x"29",x"55",x"55",x"5C",x"5D",x"35",x"27",x"27",x"56",x"4D",x"5D",x"DD",x"DC",x"18",x"C4",x"5D",x"62",x"4D",x"F3",x"63",x"B0",x"08",x"8E",x"26",x"2D",x"08",x"49",x"53",x"2D",x"5B",x"B7",x"28",x"05",x"D1",x"F0",x"5C",x"6C",x"CA",x"E0",x"24",x"D2",x"23",x"12",x"04",x"37",x"1A",x"B5",x"70",x"6B",x"AB",x"FC",x"E8",x"CD",x"43",x"BC",x"0D",x"0B",x"52",x"96",x"30",x"F3",x"A6",x"0A",x"28",x"D7",x"4C",x"03",x"21",x"CB",x"4D",x"D5",x"C4",x"5A",x"97",x"DC",x"17",x"77",x"57",x"6F",x"DC",x"2A",x"1F",x"62",x"84",x"BD",x"6D",x"AB",x"5C",x"C8",x"51",x"F2",x"AE",x"A5",x"D6",x"29",x"87",x"29",x"DA",x"B4",x"46",x"96",x"6C",x"D3",x"B4",x"DA",x"6A",x"9D",x"AA",x"1D",x"63",x"69",x"6B",x"7C",x"AC",x"31",x"CA",x"B6",x"AD",x"8D",x"A1",x"46",x"39",x"BB",x"B4",x"3E",x"B9",x"1C",x"93",x"6C",x"D3",x"86",x"E4",x"AA",x"93",x"63",x"69",x"1A",x"93",x"E9",x"2C",x"D5",x"67",x"0C",x"F0",x"2E",x"D2",x"35",x"3E",x"D4",x"18",x"45",x"9B",x"D6",x"66",x"E7",x"ED",x"EE",x"49",x"4B",x"17",x"5C",x"94",x"58",x"45",x"6A",x"43",x"2C",x"61",x"E2",x"65",x"B6",x"8D",x"B1",x"A4",x"AA",x"65",x"D1",x"30",x"FA",x"49",x"5A",x"65",x"76",x"C3",x"18",x"0E",x"6A",x"A7",x"3A",x"0B",x"63",x"3C",x"A8",x"15",x"E6",x"2C",x"8D",x"69",x"42",x"A6",x"7A",x"D6",x"36",x"A5",x"2A",x"21",x"E9",x"5D",x"DA",x"9C",x"93",x"2B",x"47",x"B7",x"1D",x"4B",x"0D",x"EE",x"E4",x"BE",x"66",x"6C",x"DD",x"85",x"B1",x"F9",x"93",x"31",x"0E",x"EB",x"C6",x"EA",x"73",x"C6",x"D8",x"AD",x"2B",x"AB",x"47",x"2D",x"63",x"F5",x"E6",x"9C",x"E6",x"BC",x"F5",x"33",x"68",x"B8",x"68",x"33",x"05",x"AC",x"96",x"D6",x"B6",x"59",x"CB",x"55",x"D8",x"5D",x"DB",x"56",x"2D",x"33",x"95",x"B8",x"65",x"9F",x"25",x"4C",x"D8",x"92",x"A6",x"35",x"29",x"49",x"99",x"58",x"DC",x"A6",x"E6",x"AC",x"C0",x"6D",x"6D",x"5B",x"8A",x"F3",x"44",x"EF",x"D6",x"65",x"AA",x"D6",x"43",x"34",x"5A",x"A7",x"75",x"38",x"15",x"13",x"4D",x"EA",x"B6",x"6E",x"49",x"D4",x"32",x"8E",x"D9",x"93",x"90",x"F0",x"CA",x"44",x"6A",x"4F",x"5A",x"53",x"32",x"12",x"B1",x"33",x"3A",x"4B",x"4A",x"8F",x"F5",x"00",x"FF",
		x"60",x"A9",x"08",x"2D",x"8B",x"B2",x"6B",x"B5",x"24",x"C5",x"2A",x"93",x"9A",x"33",x"A2",x"1C",x"32",x"CD",x"6A",x"F6",x"88",x"72",x"70",x"F3",x"E8",x"C5",x"23",x"2C",x"41",x"CC",x"BD",x"66",x"B7",x"20",x"39",x"8E",x"CC",x"9C",x"14",x"D2",x"A2",x"DC",x"DD",x"D5",x"76",x"4A",x"B3",x"CD",x"72",x"D7",x"38",x"25",x"CE",x"3E",x"D2",x"2C",x"2B",x"25",x"2F",x"7B",x"73",x"D5",x"2A",x"31",x"DC",x"EC",x"4D",x"D5",x"73",x"F2",x"70",x"92",x"D7",x"34",x"EF",x"2A",x"C3",x"CB",x"29",x"DD",x"22",x"2A",x"8F",x"20",x"E7",x"74",x"8F",x"98",x"3D",x"82",x"5C",x"CC",x"D5",x"BB",x"0A",x"10",x"80",x"47",x"0B",x"E3",x"64",x"67",x"E1",x"56",x"95",x"83",x"57",x"55",x"87",x"7B",x"C4",x"09",x"7E",x"55",x"EB",x"61",x"DE",x"5A",x"00",x"49",x"2D",x"33",x"60",x"B2",x"30",x"06",x"6C",x"1E",x"CE",x"80",x"2D",x"C3",x"18",x"B0",x"55",x"5A",x"31",x"9A",x"67",x"51",x"9D",x"CA",x"CD",x"A8",x"52",x"A4",x"7A",x"02",x"15",x"AB",x"30",x"D1",x"9E",x"36",x"5C",x"EC",x"8C",x"35",x"7A",x"42",x"48",x"71",x"0A",x"51",x"ED",x"73",x"2A",x"C5",x"AD",x"58",x"34",x"2F",x"A4",x"16",x"AF",x"63",x"91",x"58",x"93",x"DB",x"FC",x"21",x"95",x"62",x"4C",x"4E",x"09",x"9A",x"62",x"E9",x"36",x"3B",x"29",x"4A",x"4A",x"3D",x"CD",x"63",x"BB",x"38",x"28",x"8D",x"F2",x"A8",x"14",x"92",x"A0",x"DC",x"C2",x"B3",x"52",x"48",x"83",x"B4",x"48",x"8B",x"CA",x"21",x"8B",x"5C",x"62",x"5C",x"6B",x"87",x"22",x"71",x"B1",x"0A",x"6D",x"1C",x"DA",x"49",x"DC",x"49",x"3C",x"B5",x"00",x"1A",x"34",x"13",x"40",x"85",x"AE",x"0C",x"28",x"50",x"CD",x"C5",x"9D",x"B9",x"B8",x"49",x"ED",x"52",x"86",x"6C",x"6E",x"31",x"51",x"5A",x"9D",x"75",x"65",x"A8",x"DF",x"19",x"4D",x"32",x"E5",x"EE",x"79",x"7B",x"34",x"45",x"85",x"B9",x"D5",x"12",x"53",x"77",x"6D",x"AE",x"62",x"49",x"08",x"50",x"A1",x"84",x"02",x"0A",x"B5",x"72",x"40",x"53",x"1A",x"0C",x"48",x"36",x"9D",x"00",x"45",x"85",x"81",x"A9",x"BD",x"D3",x"70",x"57",x"27",x"A6",x"76",x"C3",x"C4",x"DD",x"9C",x"98",x"C6",x"1F",x"B4",x"6E",x"53",x"EB",x"EA",x"B0",x"21",x"DB",x"25",x"6B",x"AA",x"E3",x"C4",x"4C",x"93",x"AC",x"AD",x"89",x"49",x"3D",x"2D",x"96",x"8E",x"36",x"3B",x"D3",x"88",x"58",x"32",x"EA",x"62",x"4D",x"AD",x"6A",x"C9",x"E8",x"AB",x"35",x"E5",x"CA",x"37",x"A3",x"EF",x"36",x"94",x"C2",x"D7",x"94",x"AE",x"24",x"36",x"4B",x"69",x"EC",x"9A",x"94",x"CC",x"DC",x"3D",x"6D",x"68",x"B3",x"37",x"0D",x"8B",x"CA",x"A9",x"8F",x"DE",x"D4",x"DC",x"ED",x"B6",x"3E",x"5A",x"77",x"4D",x"8B",x"DB",x"FA",x"E8",x"C2",x"34",x"2D",x"6E",x"E8",x"43",x"23",x"CF",x"B4",x"C4",x"A1",x"8F",x"0D",x"23",x"4B",x"B2",x"A4",x"21",x"55",x"8C",x"4C",x"EB",x"DC",x"C6",x"9C",x"44",x"2D",x"7D",x"CD",x"98",x"AA",x"35",x"95",x"88",x"25",x"63",x"6A",x"D6",x"95",x"BD",x"96",x"8C",x"A9",x"1B",x"33",x"8A",x"5C",x"D2",x"E6",x"AE",x"4D",x"29",x"72",x"49",x"99",x"87",x"54",x"95",x"C8",x"25",x"65",x"E9",x"4A",x"45",x"B2",x"E6",x"86",x"AD",x"3A",x"11",x"EE",x"A8",x"A7",x"F6",x"68",x"CD",x"AC",x"23",x"2A",x"3B",x"83",x"D2",x"88",x"71",x"43",x"0F",x"FF",
		x"60",x"A2",x"8C",x"CA",x"D4",x"C3",x"6C",x"A7",x"3C",x"5A",x"73",x"AB",x"AA",x"3C",x"F2",x"EC",x"2D",x"A4",x"EA",x"F2",x"28",x"8B",x"F7",x"94",x"CA",x"2B",x"23",x"2F",x"21",x"8A",x"2B",x"6F",x"8F",x"24",x"FB",x"4C",x"AD",x"6A",x"34",x"FC",x"18",x"43",x"BB",x"DB",x"CE",x"F0",x"8B",x"37",x"53",x"5F",x"27",x"C0",x"80",x"EC",x"34",x"52",x"59",x"BC",x"A7",x"54",x"5E",x"49",x"71",x"F1",x"51",x"5C",x"71",x"B9",x"C4",x"D9",x"47",x"70",x"45",x"C8",x"94",x"F8",x"18",x"56",x"1E",x"52",x"5A",x"16",x"92",x"97",x"A8",x"67",x"1E",x"79",x"48",x"96",x"66",x"B5",x"78",x"94",x"C1",x"87",x"66",x"56",x"E3",x"D6",x"14",x"E3",x"2E",x"1C",x"9B",x"04",x"10",x"51",x"88",x"00",x"22",x"2E",x"6D",x"55",x"F2",x"6E",x"AA",x"5D",x"7B",x"D4",x"29",x"86",x"89",x"77",x"E3",x"D1",x"26",x"1F",x"61",x"56",x"6D",x"46",x"9F",x"B2",x"27",x"57",x"36",x"6A",x"63",x"B6",x"5E",x"6E",x"11",x"B3",x"75",x"29",x"66",x"86",x"46",x"AC",x"D6",x"A6",x"1C",x"69",x"92",x"B6",x"5A",x"1D",x"9B",x"15",x"7B",x"36",x"6A",x"75",x"C8",x"9A",x"E6",x"DE",x"B9",x"D5",x"BE",x"A8",x"7B",x"86",x"D7",x"54",x"87",x"2A",x"21",x"E1",x"4A",x"53",x"15",x"06",x"B9",x"BB",x"7A",x"2B",x"55",x"C8",x"94",x"2D",x"D1",x"76",x"D4",x"31",x"59",x"9A",x"65",x"9B",x"D1",x"44",x"9B",x"19",x"62",x"4B",x"47",x"1B",x"6D",x"74",x"88",x"AD",x"19",x"5D",x"70",x"D1",x"C1",x"B6",x"75",x"74",x"C9",x"66",x"06",x"4B",x"B7",x"D1",x"25",x"17",x"69",x"AC",x"5B",x"47",x"9F",x"BD",x"87",x"99",x"6D",x"1E",x"43",x"B1",x"6A",x"9A",x"DA",x"39",x"35",x"C9",x"7A",x"94",x"EA",x"52",x"D6",x"46",x"17",x"1D",x"E2",x"5B",x"04",x"90",x"AC",x"26",x"05",x"CA",x"94",x"83",x"BA",x"4D",x"4D",x"19",x"5D",x"0D",x"1E",x"92",x"7E",x"65",x"74",x"25",x"5A",x"72",x"C5",x"94",x"31",x"94",x"6C",x"29",x"16",x"8D",x"43",x"9F",x"AD",x"99",x"BB",x"37",x"66",x"40",x"91",x"AE",x"02",x"A8",x"26",x"AD",x"B4",x"B5",x"BA",x"85",x"A8",x"D3",x"D2",x"C6",x"22",x"66",x"6D",x"F5",x"4A",x"93",x"3A",x"6B",x"A4",x"35",x"2B",x"65",x"6A",x"A4",x"99",x"BE",x"26",x"25",x"B9",x"42",x"A6",x"E7",x"22",x"17",x"D7",x"28",x"AC",x"11",x"6D",x"80",x"00",x"C5",x"87",x"33",x"20",x"A8",x"52",x"04",x"F8",x"8C",x"F3",x"00",x"FF",
		x"60",x"04",x"18",x"32",x"8C",x"00",x"5B",x"3B",x"13",x"60",x"AB",x"30",x"02",x"1C",x"11",x"9A",x"86",x"26",x"45",x"9B",x"6C",x"51",x"EB",x"9A",x"95",x"16",x"D3",x"CD",x"AD",x"6D",x"4E",x"47",x"45",x"FB",x"8C",x"A6",x"19",x"99",x"10",x"EB",x"3A",x"EA",x"AA",x"6C",x"92",x"B5",x"6D",x"AB",x"B3",x"C8",x"0C",x"E2",x"26",x"A5",x"CA",x"8C",x"6D",x"4D",x"E3",x"96",x"2A",x"51",x"B6",x"33",x"89",x"DB",x"EA",x"28",x"3D",x"83",x"2C",x"72",x"6B",x"A2",x"B6",x"31",x"89",x"9A",x"AD",x"8D",x"2A",x"37",x"D8",x"12",x"B7",x"2E",x"89",x"9C",x"22",x"59",x"DA",x"FA",x"2C",x"63",x"92",x"74",x"ED",x"E8",x"AB",x"88",x"74",x"F5",x"D6",x"63",x"68",x"32",x"83",x"CD",x"5B",x"95",x"A1",x"28",x"0E",x"E7",x"A8",x"52",x"86",x"A2",x"24",x"43",x"A3",x"4C",x"E9",x"B3",x"F0",x"0A",x"B5",x"C8",x"65",x"28",x"52",x"AB",x"58",x"1D",x"97",x"A9",x"C8",x"A8",x"20",x"69",x"5C",x"86",x"C2",x"3D",x"4D",x"BC",x"56",x"E8",x"A7",x"D1",x"50",x"53",x"37",x"02",x"98",x"96",x"51",x"00",x"33",x"08",x"09",x"60",x"14",x"33",x"01",x"8C",x"26",x"DA",x"A2",x"DE",x"DC",x"54",x"24",x"59",x"4B",x"62",x"36",x"8D",x"EC",x"CA",x"2D",x"CD",x"76",x"22",x"D9",x"1F",x"B7",x"2C",x"9B",x"89",x"54",x"BF",x"DD",x"D2",x"EC",x"D7",x"C3",x"72",x"4A",x"48",x"62",x"8A",x"B4",x"98",x"28",x"0C",x"C8",x"92",x"8B",x"00",x"CD",x"A3",x"B9",x"38",x"46",x"D7",x"A8",x"AA",x"5C",x"D2",x"6C",x"3B",x"52",x"62",x"4E",x"CB",x"B2",x"99",x"48",x"B5",x"DA",x"2D",x"8A",x"D1",x"4C",x"6D",x"C7",x"B4",x"C4",x"DB",x"48",x"F7",x"68",x"64",x"8A",x"6C",x"CC",x"54",x"CD",x"2E",x"02",x"A2",x"34",x"45",x"40",x"D4",x"66",x"08",x"C8",x"DA",x"15",x"01",x"96",x"AB",x"87",x"30",x"D9",x"50",x"8B",x"6A",x"92",x"E2",x"E8",x"CD",x"CD",x"2D",x"76",x"89",x"43",x"D0",x"12",x"F1",x"55",x"2D",x"F3",x"D1",x"DD",x"B1",x"3B",x"B7",x"DC",x"B9",x"F4",x"A4",x"EA",x"DC",x"CA",x"60",x"C3",x"12",x"BD",x"6F",x"6B",x"22",x"2F",x"2B",x"32",x"7F",x"AD",x"8D",x"3A",x"3C",x"48",x"FC",x"B5",x"2E",x"8A",x"B4",x"62",x"F5",x"D7",x"FA",x"AC",x"DC",x"4B",x"44",x"5F",x"1B",x"93",x"0A",x"2F",x"66",x"FF",x"65",x"8A",x"C2",x"3D",x"55",x"F5",x"95",x"29",x"18",x"8F",x"60",x"CD",x"97",x"E6",x"A8",x"2C",x"DC",x"58",x"7F",x"59",x"A2",x"B6",x"30",x"E3",x"7C",x"65",x"C9",x"46",x"4C",x"43",x"FD",x"85",x"39",x"07",x"21",x"F3",x"B0",x"4D",x"96",x"24",x"DD",x"8A",x"45",x"AB",x"5B",x"BB",x"D5",x"92",x"70",x"C9",x"62",x"AE",x"8A",x"C3",x"CD",x"A3",x"B0",x"35",x"0B",x"75",x"77",x"57",x"F2",x"00",x"FF",
		x"60",x"89",x"EE",x"51",x"5C",x"32",x"A3",x"26",x"BA",x"F7",x"0E",x"72",x"1B",x"DB",x"E8",x"9E",x"CB",x"68",x"BC",x"72",x"62",x"9B",x"51",x"D3",x"8B",x"30",x"0C",x"48",x"8A",x"D5",x"70",x"D5",x"B1",x"79",x"59",x"94",x"45",x"AF",x"10",x"89",x"99",x"4D",x"12",x"3D",x"73",x"0D",x"6A",x"8D",x"59",x"EC",x"0A",x"9E",x"14",x"59",x"A5",x"48",x"9D",x"4B",x"78",x"A7",x"19",x"04",x"08",x"15",x"D5",x"C4",x"1E",x"45",x"B5",x"B2",x"DC",x"E2",x"7B",x"0E",x"E3",x"F4",x"C9",x"45",x"E9",x"2E",x"98",x"CE",x"42",x"13",x"C0",x"B1",x"08",x"04",x"74",x"19",x"16",x"F4",x"EE",x"5D",x"B5",x"AC",x"F2",x"90",x"5A",x"4E",x"A1",x"F2",x"29",x"43",x"6E",x"4D",x"4D",x"32",x"CA",x"26",x"AB",x"45",x"17",x"39",x"8F",x"8C",x"00",x"67",x"38",x"10",x"40",x"6D",x"66",x"B1",x"DB",x"74",x"E3",x"88",x"B1",x"C5",x"6C",x"DD",x"9C",x"3D",x"A6",x"06",x"B7",x"15",x"63",x"3D",x"8F",x"8C",x"80",x"64",x"C1",x"00",x"01",x"D6",x"5A",x"36",x"BF",x"F7",x"4E",x"0A",x"99",x"DD",x"DC",x"76",x"B3",x"D8",x"75",x"6A",x"F1",x"DA",x"F3",x"26",x"8F",x"BA",x"C3",x"6F",x"2F",x"4B",x"CC",x"AA",x"8E",x"B0",x"3D",x"4F",x"09",x"9B",x"DA",x"E2",x"FA",x"AC",x"D8",x"7C",x"6E",x"C9",x"DA",x"B6",x"62",x"B7",x"A9",x"2E",x"AF",x"DD",x"9C",x"D3",x"A7",x"3C",x"FF",
		x"60",x"CE",x"9B",x"52",x"14",x"A7",x"E2",x"34",x"AB",x"97",x"60",x"74",x"9F",x"DA",x"CC",x"F6",x"AC",x"88",x"BC",x"1E",x"73",x"B2",x"43",x"8E",x"CC",x"46",x"20",x"80",x"AA",x"35",x"92",x"5A",x"95",x"86",x"B6",x"4B",x"1E",x"CA",x"F0",x"1E",x"D8",x"1D",x"65",x"A8",x"33",x"45",x"51",x"56",x"B5",x"A1",x"8D",x"D2",x"8D",x"11",x"95",x"87",x"D6",x"4B",x"27",x"94",x"C7",x"16",x"56",x"B1",x"C4",x"3A",x"29",x"05",x"80",x"01",x"CD",x"6B",x"0A",x"60",x"58",x"89",x"A6",x"D7",x"A0",x"E6",x"AB",x"B1",x"87",x"D6",x"63",x"17",x"66",x"56",x"1D",x"5A",x"4F",x"3D",x"94",x"51",x"75",x"E8",x"33",x"46",x"63",x"66",x"DC",x"64",x"0C",x"EB",x"8E",x"15",x"B6",x"11",x"A0",x"A5",x"39",x"01",x"2A",x"0B",x"55",x"C0",x"0E",x"A9",x"0C",x"30",x"5A",x"8B",x"C9",x"D1",x"A8",x"85",x"6B",x"22",x"23",x"66",x"2B",x"E6",x"41",x"2D",x"13",x"D3",x"9D",x"AB",x"B4",x"3B",x"59",x"F4",x"C9",x"11",x"64",x"D5",x"74",x"D1",x"B7",x"B9",x"78",x"44",x"AB",x"45",x"DF",x"E6",x"E2",x"11",x"8D",x"06",x"F5",x"7A",x"8A",x"AA",x"35",x"1A",x"F4",x"4B",x"9D",x"84",x"59",x"65",x"30",x"BF",x"86",x"09",x"67",x"ED",x"C1",x"FE",x"12",x"4E",x"5C",x"55",x"07",x"FF",x"62",x"27",x"52",x"57",x"69",x"FC",x"4F",x"AE",x"A8",x"13",x"B7",x"88",x"D7",x"B0",x"48",x"95",x"12",x"23",x"37",x"A8",x"D5",x"1D",x"76",x"8D",x"DE",x"A0",x"64",x"97",x"DB",x"79",x"FF",
		x"60",x"4E",x"2D",x"9B",x"2B",x"2C",x"EB",x"14",x"BE",x"6C",x"1A",x"AB",x"4A",x"32",x"98",x"72",x"B4",x"24",x"62",x"CE",x"60",x"4B",x"D6",x"F2",x"CA",x"A8",x"49",x"CA",x"C5",x"AD",x"2A",x"CC",x"20",x"20",x"26",x"F1",x"C1",x"96",x"6A",x"2D",x"13",x"71",x"06",x"53",x"A6",x"15",x"CF",x"C4",x"1E",x"6C",x"29",x"DE",x"5C",x"93",x"7A",x"88",x"A5",x"45",x"53",x"57",x"D4",x"A2",x"A5",x"2E",x"65",x"1B",x"72",x"87",x"98",x"B7",x"A5",x"74",x"45",x"1B",x"5C",x"89",x"36",x"DC",x"93",x"64",x"08",x"A5",x"78",x"4B",x"56",x"BD",x"A1",x"A5",x"61",x"E9",x"5D",x"61",x"9D",x"93",x"BA",x"7B",x"46",x"49",x"1D",x"5A",x"EA",x"5A",x"DE",x"15",x"75",x"48",x"A5",x"FA",x"50",x"55",x"DC",x"C1",x"D7",x"64",x"4B",x"31",x"69",x"87",x"50",x"B3",x"8D",x"44",x"D6",x"1B",x"72",x"AD",x"BE",x"38",x"99",x"64",x"C8",x"A5",x"C7",x"50",x"65",x"93",x"A1",x"94",x"E2",x"8B",x"E3",x"49",x"86",x"5E",x"AA",x"0D",x"4E",x"C6",x"19",x"66",x"A9",x"36",x"78",x"99",x"A4",x"D9",x"25",x"EB",x"D0",x"65",x"93",x"E4",x"96",x"62",x"8D",x"1F",x"A9",x"BC",x"A7",x"7D",x"1C",x"3E",x"FF",
		x"60",x"C1",x"E8",x"81",x"02",x"D6",x"13",x"37",x"B5",x"76",x"4E",x"D6",x"F4",x"1D",x"B4",x"3C",x"A8",x"C1",x"3B",x"2D",x"00",x"80",x"00",x"9A",x"36",x"1D",x"7C",x"2D",x"62",x"96",x"55",x"75",x"B0",x"2D",x"99",x"69",x"FB",x"B4",x"46",x"B7",x"6E",x"26",x"93",x"75",x"0B",x"DD",x"6B",x"38",x"75",x"4C",x"0D",x"7C",x"F5",x"6A",x"D6",x"5A",x"17",x"01",x"C1",x"AA",x"03",x"01",x"5A",x"D2",x"14",x"40",x"73",x"6C",x"43",x"2E",x"5E",x"B5",x"CB",x"8B",x"2C",x"A5",x"85",x"54",x"19",x"9F",x"BD",x"D4",x"1E",x"D2",x"34",x"7C",x"9C",x"B1",x"B3",x"12",x"53",x"8F",x"20",x"40",x"80",x"2A",x"42",x"05",x"70",x"7C",x"28",x"03",x"8A",x"66",x"61",x"4A",x"97",x"61",x"6E",x"66",x"DB",x"48",x"D1",x"E3",x"B8",x"A4",x"95",x"46",x"96",x"C5",x"E1",x"1A",x"71",x"07",x"31",x"5C",x"3A",x"8D",x"4F",x"1A",x"C4",x"F1",x"9A",x"5C",x"99",x"68",x"10",x"37",x"68",x"48",x"56",x"B9",x"41",x"6E",x"3F",x"03",x"BA",x"51",x"06",x"75",x"5C",x"16",x"68",x"56",x"19",x"D4",x"F0",x"65",x"E0",x"55",x"79",x"50",x"3D",x"87",x"40",x"66",x"9C",x"41",x"F5",x"60",x"82",x"DE",x"71",x"06",x"33",x"AC",x"0B",x"65",x"44",x"1E",x"EC",x"70",x"4D",x"30",x"19",x"2B",x"88",x"4D",x"1B",x"C5",x"49",x"E4",x"07",x"FF",
		x"60",x"04",x"C8",x"9A",x"73",x"29",x"AD",x"64",x"C8",x"B8",x"ED",x"25",x"B6",x"1A",x"61",x"65",x"76",x"96",x"D8",x"4B",x"85",x"B6",x"D9",x"5E",x"72",x"CF",x"93",x"9A",x"11",x"7B",x"E9",x"23",x"75",x"58",x"59",x"E4",x"61",x"F5",x"E8",x"66",x"61",x"76",x"93",x"3D",x"A2",x"9B",x"A8",x"C7",x"66",x"40",x"D2",x"64",x"C3",x"EC",x"25",x"9D",x"CB",x"E2",x"2C",x"BD",x"E7",x"4C",x"6E",x"8F",x"B3",x"CC",x"51",x"2A",x"B9",x"22",x"EE",x"B2",x"46",x"A9",x"A4",x"8C",x"B8",x"CB",x"1E",x"A5",x"92",x"D2",x"E3",x"2E",x"7B",x"94",x"4C",x"4A",x"8F",x"BB",x"EC",x"91",x"2B",x"29",x"23",x"EE",x"B2",x"47",x"A9",x"A0",x"F4",x"38",x"CB",x"19",x"A5",x"9C",x"D3",x"63",x"0F",x"67",x"B4",x"70",x"0D",x"AF",x"92",x"DC",x"9E",x"CC",x"CC",x"DD",x"EA",x"03",x"FF",
		x"60",x"0C",x"C8",x"55",x"7D",x"08",x"A5",x"7B",x"59",x"79",x"D5",x"C1",x"95",x"16",x"65",x"6D",x"55",x"07",x"5B",x"8B",x"8F",x"A5",x"55",x"19",x"6C",x"AB",x"9E",x"9E",x"E6",x"B4",x"71",x"B5",x"45",x"44",x"AA",x"1C",x"02",x"F8",x"40",x"16",x"84",x"52",x"2C",x"2C",x"D4",x"CE",x"10",x"6B",x"B6",x"8E",x"34",x"BB",x"43",x"6C",x"D9",x"26",x"4A",x"EB",x"0C",x"A9",x"96",x"18",x"2D",x"9B",x"32",x"E4",x"D2",x"AD",x"AD",x"6C",x"F6",x"50",x"4A",x"B5",x"F6",x"B6",x"A9",x"43",x"2D",x"C5",x"DA",x"DB",x"AE",x"0E",x"B5",x"14",x"2B",x"1F",x"BB",x"32",x"94",x"52",x"3D",x"6D",x"6D",x"4E",x"52",x"4A",x"8B",x"B0",x"72",x"3B",x"0F",x"FF",
		x"60",x"08",x"28",x"5E",x"CD",x"31",x"35",x"4A",x"9B",x"7B",x"AC",x"25",x"D4",x"E4",x"A3",x"E9",x"4E",x"16",x"DF",x"B2",x"97",x"57",x"58",x"5D",x"5C",x"EB",x"5E",x"D6",x"11",x"76",x"71",x"BD",x"45",x"5B",x"5A",x"B4",x"C5",x"F5",x"9A",x"6D",x"61",x"51",x"17",x"DB",x"6A",x"25",x"A7",x"3B",x"29",x"4C",x"6D",x"19",x"96",x"26",x"27",x"D1",x"B5",x"99",x"5B",x"88",x"53",x"27",x"D7",x"66",x"2E",x"AA",x"B2",x"93",x"9C",x"AB",x"15",x"B7",x"DA",x"6A",x"4A",x"5E",x"96",x"B2",x"69",x"B9",x"A9",x"A9",x"7B",x"E9",x"74",x"E4",x"A6",x"A6",x"E1",x"A5",x"D3",x"91",x"9B",x"9A",x"BB",x"97",x"4C",x"D7",x"6E",x"6A",x"6E",x"51",x"3A",x"55",x"A7",x"A9",x"B9",x"47",x"C9",x"7A",x"DC",x"A6",x"E5",x"E9",x"A9",x"63",x"76",x"92",x"52",x"A7",x"B7",x"96",x"45",x"2A",x"62",x"AD",x"D6",x"52",x"6A",x"6B",x"F0",x"B5",x"5A",x"59",x"AB",x"93",x"C5",x"B5",x"E6",x"65",x"99",x"51",x"17",x"D7",x"AB",x"B7",x"65",x"46",x"5D",x"5C",x"6B",x"51",x"1A",x"11",x"75",x"71",x"AD",x"45",x"69",x"44",x"DC",x"C5",x"B5",x"16",x"A5",x"E1",x"76",x"17",x"57",x"9B",x"A5",x"A5",x"39",x"6D",x"7C",x"1D",x"9A",x"D1",x"A2",x"A4",x"88",x"A5",x"59",x"6B",x"89",x"CD",x"22",x"E5",x"69",x"49",x"6D",x"96",x"86",x"94",x"87",x"17",x"4F",x"58",x"1E",x"72",x"9E",x"9E",x"3A",x"65",x"B9",x"29",x"79",x"78",x"C9",x"B6",x"E5",x"A6",x"E6",x"E1",x"C5",x"DB",x"91",x"9B",x"9A",x"9B",x"37",x"4F",x"D7",x"29",x"6A",x"AE",x"D1",x"D2",x"5D",x"27",x"69",x"B9",x"7A",x"C9",x"54",x"9C",x"A0",x"97",x"65",x"21",x"ED",x"89",x"1F",x"FF",
		x"60",x"22",x"B0",x"4E",x"53",x"BA",x"6C",x"06",x"D3",x"19",x"49",x"ED",x"88",x"99",x"74",x"A7",x"B5",x"B4",x"C3",x"66",x"51",x"AC",x"B5",x"B0",x"76",x"9B",x"45",x"0E",x"4E",x"5D",x"27",x"14",x"16",x"39",x"38",x"0E",x"CF",x"70",x"D0",x"E4",x"18",x"D8",x"34",x"B3",x"56",x"93",x"83",x"67",x"B3",x"8A",x"58",x"C9",x"10",x"DA",x"3D",x"32",x"12",x"39",x"DF",x"73",x"77",x"8F",x"88",x"65",x"8A",x"24",x"58",x"23",x"33",x"B5",x"4A",x"02",x"57",x"0D",x"8F",x"34",x"C6",x"17",x"4E",x"DC",x"23",x"23",x"05",x"CB",x"04",x"36",x"8F",x"B4",x"9D",x"74",x"ED",x"39",x"22",x"C3",x"51",x"50",x"4D",x"10",x"B7",x"8E",x"58",x"49",x"B5",x"91",x"DD",x"2A",x"62",x"05",x"D5",x"44",x"F6",x"C8",x"B0",x"15",x"34",x"9B",x"D8",x"3D",x"CC",x"76",x"D2",x"75",x"50",x"77",x"77",x"39",x"49",x"37",x"C1",x"DC",x"42",x"94",x"04",x"43",x"47",x"71",x"4B",x"51",x"E2",x"4C",x"19",x"D4",x"AC",x"43",x"96",x"B1",x"A9",x"8B",x"88",x"4C",x"47",x"C6",x"E5",x"DA",x"2C",x"B3",x"12",x"2B",x"DF",x"6B",x"61",x"CD",x"4C",x"23",x"22",x"2F",x"4C",x"3C",x"32",x"31",x"C9",x"BB",x"0C",x"73",x"33",x"DB",x"0F",x"FF",
		x"60",x"08",x"F0",x"0E",x"4D",x"89",x"C9",x"51",x"64",x"46",x"4C",x"63",x"C7",x"C4",x"1D",x"55",x"96",x"93",x"1A",x"13",x"67",x"B6",x"85",x"49",x"A2",x"8F",x"32",x"3E",x"19",x"B6",x"88",x"BE",x"C8",x"64",x"A6",x"95",x"22",x"86",x"C4",x"1D",x"55",x"96",x"93",x"18",x"32",x"4D",x"74",x"45",x"4E",x"82",x"AF",x"BC",x"95",x"11",x"37",x"09",x"21",x"D3",x"44",x"45",x"D8",x"26",x"E5",x"4C",x"69",x"15",x"65",x"8A",x"94",x"32",x"55",x"94",x"87",x"49",x"B2",x"4F",x"3C",x"6E",x"11",x"BB",x"28",x"A9",x"60",x"59",x"7B",x"94",x"A2",x"E5",x"46",x"21",x"61",x"55",x"92",x"91",x"0B",x"26",x"87",x"47",x"4E",x"76",x"29",x"94",x"1C",x"1E",x"29",x"B8",x"29",x"52",x"5B",x"79",x"C5",x"10",x"E4",x"46",x"21",x"11",x"16",x"4D",x"92",x"2B",x"BB",x"A6",x"5B",x"74",x"79",x"1D",x"6A",x"94",x"6A",x"D3",x"15",x"25",x"AB",x"4B",x"69",x"4C",x"56",x"D6",x"22",x"CA",x"AE",x"11",x"1E",x"FF",
		x"60",x"46",x"63",x"21",x"3C",x"C3",x"2D",x"3B",x"39",x"04",x"71",x"CB",x"90",x"EC",x"B8",x"98",x"25",x"B8",x"5D",x"66",x"92",x"B4",x"D7",x"D4",x"76",x"39",x"49",x"36",x"5E",x"DD",x"D2",x"E4",x"04",x"5E",x"25",x"0D",x"5D",x"55",x"EC",x"38",x"5F",x"35",x"25",x"D9",x"49",x"92",x"B5",x"D7",x"B4",x"0C",x"59",x"C9",x"30",x"4E",x"DC",x"32",x"6C",x"07",x"43",x"79",x"C9",x"08",x"53",x"E2",x"2C",x"6D",x"C5",x"BD",x"C2",x"B6",x"73",x"9D",x"61",x"97",x"4E",x"C5",x"CA",x"F7",x"46",x"4C",x"B2",x"1C",x"89",x"38",x"08",x"56",x"0B",x"4B",x"CC",x"B2",x"24",x"54",x"CC",x"3D",x"31",x"8B",x"3D",x"57",x"B1",x"F0",x"D8",x"2C",x"0E",x"4A",x"45",x"3D",x"12",x"B3",x"BC",x"CB",x"30",x"37",x"B3",x"FD",x"00",x"FF",
		x"60",x"42",x"CD",x"19",x"9D",x"D3",x"13",x"05",x"D5",x"27",x"EE",x"18",x"B1",x"58",x"54",x"9F",x"68",x"A3",x"D2",x"52",x"53",x"43",x"A4",x"89",x"CE",x"98",x"4D",x"CF",x"09",x"53",x"DB",x"2B",x"36",x"23",x"67",x"2C",x"6D",x"0F",x"D5",x"EC",x"94",x"A8",x"B4",x"AD",x"70",x"73",x"53",x"A6",x"F4",x"D1",x"D0",x"C5",x"CB",x"95",x"42",x"4B",x"87",x"94",x"20",x"15",x"2A",x"2B",x"AD",x"9C",x"E2",x"50",x"B8",x"DC",x"DD",x"52",x"48",x"53",x"A4",x"4A",x"73",x"53",x"21",x"CB",x"19",x"D3",x"2C",x"2C",x"B9",x"BC",x"34",x"74",x"F6",x"B4",x"E8",x"AA",x"3A",x"C9",x"89",x"C3",x"96",x"A9",x"CB",x"64",x"13",x"31",x"5B",x"A2",x"2E",x"9D",x"5D",x"D8",x"2C",x"3D",x"FF",
		x"60",x"CA",x"8A",x"5E",x"25",x"2C",x"A7",x"38",x"4B",x"55",x"A9",x"A9",x"8E",x"9C",x"14",x"1F",x"B5",x"C2",x"BB",x"64",x"92",x"5C",x"B0",x"4E",x"CD",x"8A",x"49",x"B4",x"D9",x"32",x"D4",x"6A",x"25",x"C1",x"37",x"75",x"D7",x"58",x"94",x"C4",x"B0",x"54",x"4D",x"73",x"51",x"12",x"5D",x"77",x"31",x"8F",x"99",x"49",x"34",x"C5",x"CD",x"C5",x"6B",x"27",x"49",x"E6",x"70",x"57",x"A9",x"9C",x"14",x"13",x"B2",x"DA",x"70",x"72",x"30",x"54",x"F1",x"72",x"B6",x"CB",x"C6",x"D3",x"3A",x"C3",x"8C",x"62",x"BB",x"C0",x"16",x"2B",x"C5",x"68",x"63",x"12",x"B5",x"5C",x"CD",x"72",x"B5",x"A9",x"6C",x"B3",x"34",x"F2",x"45",x"6A",x"08",x"C6",x"23",x"45",x"DC",x"3C",x"FF",
		x"60",x"C1",x"4D",x"53",x"22",x"D2",x"CB",x"14",x"2D",x"0D",x"49",x"4B",x"2F",x"1B",x"94",x"D0",x"35",x"2C",x"35",x"72",x"90",x"43",x"D5",x"34",x"77",x"53",x"41",x"F2",x"4D",x"43",x"33",x"4D",x"07",x"D9",x"6C",x"F6",x"C8",x"8C",x"9A",x"34",x"D7",x"AC",x"28",x"2B",x"4E",x"F2",x"42",x"B1",x"24",x"AB",x"4A",x"29",x"0F",x"D9",x"53",x"D8",x"17",x"84",x"D6",x"07",x"4F",x"53",x"AD",x"E5",x"86",x"E8",x"34",x"93",x"BC",x"A1",x"5A",x"42",x"8E",x"08",x"B1",x"58",x"0F",x"FF",
		x"60",x"C1",x"8F",x"4D",x"D3",x"3A",x"85",x"05",x"37",x"0C",x"C9",x"28",x"97",x"9A",x"94",x"34",x"25",x"A2",x"CA",x"58",x"51",x"D3",x"94",x"88",x"F6",x"70",x"45",x"8D",x"53",x"C3",x"DB",x"CD",x"35",x"35",x"76",x"4B",x"E9",x"92",x"D6",x"F4",x"38",x"24",x"AD",x"D2",x"6A",x"B1",x"42",x"D7",x"B2",x"4A",x"73",x"C5",x"8F",x"53",x"DD",x"33",x"8D",x"A5",x"38",x"4C",x"33",x"CF",x"0A",x"16",x"F2",x"90",x"22",x"DD",x"3D",x"68",x"68",x"52",x"B4",x"12",x"F1",x"22",x"A1",x"4F",x"D9",x"4A",x"2D",x"82",x"86",x"3E",x"25",x"4F",x"D1",x"08",x"92",x"A6",x"54",x"D2",x"CD",x"23",x"68",x"58",x"73",x"8E",x"54",x"8F",x"30",x"6A",x"49",x"A9",x"D2",x"3C",x"82",x"3E",x"FF",
		x"60",x"CE",x"4F",x"19",x"4A",x"BB",x"12",x"14",x"27",x"7A",x"6E",x"4B",x"B7",x"59",x"EC",x"E0",x"A4",x"B5",x"CD",x"66",x"72",x"A3",x"A5",x"D2",x"35",x"4B",x"29",x"88",x"8E",x"52",x"57",x"63",x"86",x"24",x"79",x"4C",x"EB",x"48",x"19",x"8A",x"E0",x"A9",x"BC",x"C3",x"66",x"A8",x"93",x"C3",x"F2",x"2A",x"8B",x"A1",x"2D",x"85",x"89",x"3D",x"EB",x"84",x"7E",x"A4",x"50",x"26",x"71",x"9C",x"BA",x"D1",x"DD",x"98",x"45",x"76",x"68",x"46",x"75",x"15",x"56",x"3B",x"A1",x"AA",x"89",x"85",x"2C",x"D2",x"98",x"3C",x"39",x"C8",x"A8",x"B6",x"15",x"B2",x"68",x"B0",x"6D",x"23",x"62",x"8A",x"82",x"E1",x"F6",x"35",x"5B",x"21",x"48",x"1E",x"DA",x"C6",x"1B",x"85",x"B0",x"44",x"28",x"99",x"4C",x"14",x"D2",x"52",x"C1",x"B9",x"23",x"51",x"28",x"72",x"82",x"F0",x"4A",x"47",x"A1",x"CA",x"01",x"C3",x"32",x"63",x"B9",x"AA",x"04",x"34",x"F1",x"4E",x"A4",x"9A",x"56",x"94",x"59",x"34",x"0D",x"02",x"BC",x"44",x"7D",x"FF",
		x"60",x"CC",x"31",x"CA",x"D4",x"23",x"E3",x"04",x"4F",x"3A",x"75",x"CF",x"94",x"E3",x"7C",x"65",x"C5",x"AD",x"4A",x"8E",x"8B",x"BC",x"12",x"D3",x"6C",x"39",x"26",x"55",x"DA",x"35",x"2A",x"63",x"BB",x"C4",x"39",x"31",x"CD",x"94",x"53",x"82",x"E0",x"C4",x"A5",x"5D",x"4E",x"F1",x"A2",x"17",x"E3",x"36",x"27",x"C5",x"8F",x"41",x"94",x"CB",x"92",x"94",x"20",x"3A",x"51",x"69",x"8B",x"5B",x"E2",x"E4",x"C5",x"B8",x"24",x"4E",x"CA",x"63",x"44",x"D7",x"D4",x"DA",x"A1",x"0A",x"11",x"DD",x"22",x"12",x"85",x"3A",x"44",x"74",x"8D",x"48",x"14",x"BA",x"98",x"30",x"D4",x"32",x"56",x"18",x"42",x"40",x"77",x"AB",x"C4",x"61",x"0A",x"81",x"5C",x"33",x"1A",x"85",x"29",x"78",x"72",x"8B",x"6C",x"14",x"46",x"1F",x"C4",x"BC",x"DC",x"51",x"E8",x"93",x"C3",x"F4",x"F4",x"98",x"AE",x"4C",x"16",x"22",x"3A",x"22",x"86",x"38",x"5A",x"EA",x"4C",x"B3",x"94",x"A2",x"E8",x"A8",x"AB",x"CD",x"72",x"09",x"A3",x"A3",x"AE",x"74",x"D3",x"29",x"8C",x"8E",x"26",x"D3",x"43",x"A7",x"28",x"7A",x"EA",x"48",x"0F",x"9D",x"E2",x"E4",x"B1",x"B5",x"C2",x"74",x"CA",x"52",x"C0",x"F6",x"72",x"53",x"21",x"4F",x"1E",x"33",x"DD",x"43",x"A6",x"B2",x"44",x"4C",x"F7",x"34",x"15",x"EA",x"E4",x"B0",x"23",x"2C",x"A4",x"6B",x"73",x"80",x"F6",x"0C",x"93",x"61",x"48",x"1E",x"2B",x"CA",x"6D",x"84",x"B9",x"64",x"08",x"AF",x"4C",x"E0",x"96",x"DA",x"45",x"59",x"2D",x"89",x"5B",x"EA",x"50",x"63",x"D3",x"B4",x"66",x"AA",x"37",x"9D",x"8D",x"1C",x"8B",x"B1",x"4D",x"55",x"31",x"8D",x"4D",x"86",x"5A",x"88",x"39",x"C2",x"E1",x"03",x"FF",
		x"60",x"86",x"0D",x"CE",x"C5",x"33",x"63",x"15",x"2E",x"44",x"CE",x"CC",x"8C",x"D4",x"A4",x"10",x"79",x"34",x"2D",x"52",x"53",x"43",x"A4",x"B6",x"4E",x"53",x"25",x"2A",x"15",x"93",x"2B",x"5B",x"96",x"B2",x"54",x"48",x"A9",x"4C",x"98",x"86",x"9A",x"C1",x"B5",x"33",x"51",x"1A",x"EA",x"04",x"A7",x"8C",x"96",x"69",x"CC",x"05",x"83",x"22",x"1B",x"85",x"25",x"27",x"56",x"76",x"6D",x"63",x"D6",x"EA",x"9D",x"59",x"DD",x"49",x"18",x"EB",x"10",x"15",x"B1",x"B4",x"A1",x"2A",x"1E",x"4D",x"DA",x"2B",x"85",x"A2",x"38",x"74",x"A9",x"88",x"6C",x"BA",x"96",x"48",x"51",x"2A",x"16",x"02",x"A2",x"46",x"43",x"40",x"59",x"24",x"04",x"28",x"C7",x"CD",x"24",x"D1",x"93",x"BA",x"79",x"E3",x"10",x"84",x"88",x"1D",x"1D",x"36",x"8B",x"97",x"3C",x"A5",x"6C",x"58",x"4A",x"6E",x"F4",x"58",x"31",x"69",x"2B",x"19",x"21",x"60",x"C7",x"B8",x"CD",x"A4",x"07",x"47",x"1D",x"9D",x"B2",x"92",x"9A",x"13",x"94",x"4F",x"5A",x"76",x"4A",x"08",x"18",x"DE",x"61",x"89",x"69",x"CE",x"93",x"67",x"76",x"A4",x"07",x"FF",
		x"60",x"A1",x"2E",x"91",x"34",x"46",x"22",x"95",x"B2",x"64",x"0C",x"4F",x"2F",x"99",x"B2",x"14",x"68",x"3C",x"2C",x"72",x"C9",x"53",x"E4",x"8E",x"B0",x"CA",x"AD",x"48",x"99",x"3B",x"D2",x"CA",x"94",x"3C",x"25",x"EE",x"08",x"AF",x"54",x"92",x"98",x"B8",x"3C",x"3D",x"56",x"09",x"62",x"E4",x"B2",x"B4",x"CA",x"29",x"08",x"89",x"D3",x"CA",x"6A",x"87",x"30",x"25",x"2C",x"AD",x"8C",x"E9",x"C2",x"18",x"31",x"3D",x"33",x"A6",x"48",x"B8",x"2E",x"8B",x"70",x"CB",x"2C",x"D5",x"DC",x"3C",x"2C",x"62",x"89",x"90",x"AB",x"88",x"32",x"8B",x"A4",x"7C",x"16",x"D3",x"DD",x"C3",x"B4",x"71",x"99",x"4F",x"8F",x"08",x"4B",x"C6",x"A5",x"36",x"23",x"3C",x"2C",x"29",x"DF",x"19",x"D1",x"88",x"B0",x"AC",x"E2",x"E2",x"51",x"C4",x"32",x"09",x"4B",x"B2",x"41",x"76",x"CF",x"C4",x"C6",x"4D",x"0E",x"32",x"AA",x"2C",x"3A",x"3B",x"3A",x"C8",x"EC",x"B0",x"E9",x"9C",x"E8",x"20",x"B3",x"C3",x"96",x"F1",x"5B",x"57",x"21",x"D6",x"24",x"04",x"A8",x"9E",x"18",x"01",x"35",x"92",x"98",x"3C",x"3A",x"8C",x"8A",x"AA",x"E4",x"F2",x"10",x"B0",x"3A",x"AB",x"B2",x"CB",x"AD",x"E7",x"EE",x"0A",x"5B",x"AA",x"4C",x"01",x"32",x"63",x"62",x"8A",x"A6",x"75",x"51",x"36",x"57",x"F2",x"00",x"FF",
		x"60",x"8C",x"2F",x"56",x"D9",x"3C",x"12",x"17",x"31",x"65",x"2C",x"AD",x"B0",x"D5",x"C4",x"9C",x"29",x"65",x"34",x"76",x"53",x"52",x"E2",x"D0",x"D1",x"D0",x"C5",x"4A",x"05",x"CB",x"DB",x"0D",x"17",x"3F",x"57",x"2C",x"DE",x"88",x"DC",x"92",x"5C",x"39",x"39",x"63",x"56",x"CB",x"63",x"A6",x"D2",x"AC",x"9A",x"A5",x"88",x"05",x"CB",x"63",x"6A",x"95",x"32",x"55",x"28",x"CB",x"6A",x"54",x"EA",x"5C",x"A0",x"79",x"2A",x"76",x"EA",x"52",x"C4",x"B2",x"D5",x"9A",x"A9",x"4F",x"11",x"DA",x"3B",x"62",x"A6",x"31",x"27",x"C8",x"A8",x"8C",x"99",x"A6",x"92",x"20",x"75",x"32",x"56",x"58",x"4B",x"06",x"8F",x"8A",x"DA",x"08",x"08",x"06",x"8C",x"00",x"3D",x"91",x"10",x"A0",x"3B",x"14",x"D3",x"64",x"83",x"E1",x"9B",x"11",x"5D",x"1D",x"35",x"65",x"8D",x"5B",x"72",x"79",x"32",x"14",x"59",x"69",x"C9",x"C5",x"C9",x"62",x"65",x"A7",x"A9",x"E0",x"47",x"4D",x"93",x"6D",x"96",x"83",x"EB",x"1D",x"4F",x"95",x"C6",x"4E",x"B6",x"73",x"D6",x"D5",x"22",x"3B",x"58",x"D9",x"42",x"E5",x"A4",x"28",x"E7",x"66",x"07",x"EE",x"5D",x"91",x"4C",x"50",x"1C",x"84",x"75",x"54",x"74",x"61",x"49",x"60",x"D6",x"11",x"DB",x"A4",x"35",x"81",x"4A",x"66",x"2C",x"93",x"17",x"87",x"CA",x"66",x"B1",x"59",x"DB",x"8C",x"2A",x"AB",x"46",x"7E",x"FF",
		x"60",x"08",x"28",x"55",x"D9",x"71",x"BE",x"6A",x"56",x"47",x"C9",x"40",x"87",x"A2",x"9D",x"E5",x"05",x"03",x"1D",x"8A",x"74",x"A5",x"1A",x"2A",x"74",x"4A",x"12",x"D1",x"3E",x"B0",x"30",x"A9",x"50",x"E4",x"64",x"A9",x"C2",x"86",x"22",x"59",x"63",x"A5",x"0A",x"17",x"B2",x"B4",x"75",x"96",x"69",x"42",x"0C",x"1A",x"D1",x"5E",x"BA",x"28",x"A9",x"88",x"69",x"58",x"E9",x"60",x"C4",x"68",x"E2",x"C5",x"85",x"9D",x"1B",x"83",x"9A",x"97",x"86",x"32",x"51",x"2E",x"66",x"E2",x"52",x"4B",x"E4",x"C5",x"85",x"61",x"99",x"E5",x"07",x"FF",
		x"60",x"06",x"CB",x"86",x"32",x"27",x"9C",x"14",x"B4",x"66",x"F4",x"0A",x"4F",x"53",x"90",x"6C",x"71",x"B2",x"AC",x"49",x"C2",x"92",x"D2",x"CC",x"12",x"6B",x"8E",x"48",x"9A",x"AA",x"5A",x"ED",x"26",x"34",x"0A",x"CF",x"58",x"AB",x"97",x"10",x"6F",x"75",x"A7",x"23",x"6D",x"43",x"B2",x"A1",x"AC",x"D1",x"68",x"86",x"8A",x"9A",x"AA",x"53",x"E2",x"04",x"2C",x"59",x"AA",x"CC",x"68",x"1A",x"30",x"2F",x"6D",x"66",x"BC",x"6E",x"C1",x"B3",x"C6",x"AC",x"B1",x"B8",x"8C",x"49",x"92",x"7D",x"96",x"E5",x"28",x"D2",x"C9",x"A8",x"1E",x"8D",x"6B",x"88",x"60",x"78",x"AE",x"B5",x"89",x"A2",x"94",x"E8",x"C9",x"D5",x"24",x"82",x"B1",x"4A",x"6B",x"57",x"13",x"33",x"D6",x"F0",x"A8",x"7E",x"57",x"4D",x"78",x"29",x"AA",x"7A",x"D2",x"31",x"11",x"0D",x"CB",x"EA",x"4E",x"27",x"0F",x"FF",
		x"60",x"C2",x"73",x"C6",x"D2",x"34",x"22",x"19",x"D9",x"19",x"69",x"B6",x"8C",x"6D",x"28",x"5D",x"C4",x"BD",x"CA",x"92",x"C3",x"93",x"A3",x"21",x"8F",x"A6",x"0E",x"4D",x"59",x"13",x"C3",x"36",x"39",x"38",x"79",x"1E",x"4A",x"4F",x"A4",x"A0",x"14",x"75",x"24",x"29",x"BD",x"01",x"53",x"B4",x"16",x"E7",x"74",x"06",x"4C",x"25",x"4A",x"42",x"E2",x"19",x"30",x"15",x"2F",x"75",x"49",x"6A",x"C0",x"9C",x"64",x"42",x"A9",x"4D",x"80",x"8A",x"D5",x"96",x"A6",x"B8",x"01",x"CE",x"46",x"87",x"C3",x"5D",x"05",x"24",x"45",x"69",x"91",x"4A",x"14",x"B0",x"18",x"AD",x"21",x"3A",x"B2",x"23",x"7C",x"D2",x"A2",x"6C",x"B9",x"86",x"56",x"C5",x"C3",x"2C",x"2D",x"2B",x"96",x"D7",x"48",x"D3",x"B4",x"AC",x"24",x"99",x"DC",x"D5",x"CA",x"92",x"D2",x"74",x"52",x"55",x"2F",x"DB",x"CA",x"F0",x"C1",x"4C",x"3C",x"A3",x"28",x"CB",x"25",x"13",x"89",x"B4",x"AD",x"5C",x"EF",x"CD",x"D8",x"CA",x"8E",x"F2",x"BD",x"37",x"63",x"2F",x"C7",x"2A",x"0C",x"DE",x"8D",x"AD",x"6C",x"93",x"D4",x"07",x"17",x"F3",x"B4",x"FD",x"00",x"FF",
		x"60",x"89",x"29",x"D9",x"1A",x"CB",x"63",x"15",x"A2",x"B4",x"58",x"4C",x"8F",x"59",x"B0",x"92",x"78",x"A4",x"D4",x"49",x"41",x"6B",x"E1",x"B6",x"E1",x"38",x"05",x"6D",x"95",x"5B",x"46",x"62",x"17",x"AC",x"16",x"6A",x"BD",x"90",x"DC",x"88",x"5A",x"A4",x"74",x"AC",x"71",x"A3",x"4A",x"B5",x"65",x"97",x"26",x"85",x"2D",x"49",x"97",x"DD",x"12",x"27",x"31",x"17",x"6B",x"AC",x"8C",x"15",x"B4",x"54",x"AD",x"A8",x"CA",x"B2",x"71",x"62",x"B7",x"E2",x"6A",x"CB",x"2C",x"8C",x"CD",x"C3",x"A2",x"43",x"3D",x"FF",
		x"60",x"8A",x"37",x"A5",x"2A",x"95",x"33",x"1A",x"C2",x"8E",x"76",x"65",x"C9",x"A2",x"10",x"BE",x"3B",x"22",x"22",x"B1",x"42",x"F8",x"E9",x"C8",x"8C",x"C4",x"06",x"65",x"73",x"C3",x"33",x"9C",x"08",x"9C",x"CD",x"49",x"73",x"4F",x"A3",x"28",x"36",x"C6",x"44",x"3D",x"AD",x"E2",x"E5",x"1A",x"63",x"16",x"27",x"C4",x"62",x"6D",x"D3",x"85",x"E5",x"3C",x"FF",
		x"60",x"82",x"54",x"69",x"C2",x"44",x"9D",x"18",x"DC",x"EC",x"22",x"B1",x"CC",x"62",x"10",x"B1",x"2A",x"CC",x"62",x"8B",x"81",x"C5",x"A8",x"0E",x"F1",x"2D",x"02",x"E1",x"6F",x"C2",x"3C",x"BB",x"08",x"94",x"9D",x"09",x"89",x"4A",x"23",x"70",x"36",x"C7",x"C5",x"33",x"8D",x"A0",x"58",x"9D",x"10",x"B1",x"B4",x"8C",x"17",x"6B",x"8C",x"D8",x"9C",x"30",x"8D",x"D7",x"0D",x"65",x"71",x"8A",x"1C",x"E1",x"A7",x"42",x"55",x"F6",x"03",x"FF",
		x"60",x"46",x"8C",x"23",x"DD",x"75",x"42",x"17",x"36",x"07",x"DB",x"A0",x"B6",x"93",x"C8",x"D4",x"62",x"39",x"2C",x"4E",x"C0",x"D3",x"89",x"92",x"F0",x"38",x"09",x"4B",x"23",x"46",x"C2",x"92",x"24",x"32",x"67",x"3B",x"0D",x"B7",x"9D",x"98",x"3C",x"63",x"55",x"D2",x"75",x"10",x"72",x"B7",x"C1",x"4A",x"5B",x"4E",x"4D",x"D3",x"9A",x"B3",x"2D",x"19",x"27",x"75",x"1F",x"B6",x"72",x"8C",x"80",x"78",x"38",x"1F",x"FF",
		x"60",x"81",x"0B",x"DD",x"34",x"33",x"9B",x"06",x"3C",x"9E",x"10",x"4B",x"77",x"12",x"B0",x"F4",x"53",x"28",x"DB",x"6C",x"42",x"63",x"0F",x"96",x"6E",x"61",x"01",x"8B",x"47",x"D9",x"3A",x"42",x"1B",x"DA",x"37",x"35",x"CF",x"34",x"CC",x"0C",x"EF",x"5B",x"C5",x"BD",x"D4",x"03",x"FF",
		x"60",x"8A",x"E4",x"CD",x"2D",x"B2",x"6A",x"05",x"C2",x"67",x"57",x"B1",x"6A",x"14",x"F0",x"30",x"45",x"B4",x"AA",x"B1",x"C3",x"E3",x"43",x"F6",x"AD",x"D8",x"01",x"0F",x"8B",x"49",x"AF",x"62",x"1B",x"22",x"4C",x"21",x"9D",x"AE",x"ED",x"28",x"3F",x"84",x"B4",x"A6",x"B1",x"63",x"44",x"8A",x"10",x"ED",x"26",x"8E",x"97",x"35",x"44",x"2C",x"E2",x"28",x"49",x"16",x"67",x"8B",x"B4",x"23",x"74",x"96",x"D2",x"DC",x"DD",x"36",x"73",x"99",x"2F",x"53",x"F3",x"34",x"24",x"90",x"7A",x"C2",x"D4",x"92",x"3C",x"FF",
		x"60",x"C5",x"29",x"7A",x"53",x"8A",x"B2",x"14",x"35",x"C7",x"F1",x"08",x"DA",x"54",x"F8",x"D8",x"42",x"43",x"A6",x"4A",x"A2",x"D3",x"55",x"F5",x"CE",x"C6",x"06",x"4D",x"DF",x"85",x"D7",x"AC",x"04",x"24",x"16",x"2D",x"76",x"AF",x"6C",x"E0",x"90",x"BD",x"C9",x"75",x"AE",x"81",x"7D",x"F7",x"84",x"F2",x"B5",x"06",x"31",x"23",x"9C",x"2B",x"DB",x"1A",x"44",x"CE",x"54",x"CD",x"4A",x"AA",x"70",x"33",x"D3",x"30",x"DC",x"AD",x"60",x"64",x"9F",x"10",x"71",x"C7",x"C2",x"67",x"79",x"D2",x"CC",x"63",x"B3",x"58",x"96",x"49",x"25",x"71",x"42",x"0A",x"ED",x"37",x"5C",x"CC",x"D6",x"03",x"FF",
		x"60",x"C6",x"6D",x"DC",x"D1",x"6D",x"AA",x"04",x"63",x"13",x"27",x"B4",x"9C",x"13",x"A4",x"45",x"8C",x"31",x"7B",x"8A",x"C1",x"AB",x"36",x"F2",x"1E",x"3B",x"09",x"4E",x"D2",x"BC",x"B3",x"93",x"14",x"28",x"05",x"CB",x"C8",x"4E",x"9A",x"D0",x"D4",x"BC",x"35",x"3B",x"59",x"42",x"D2",x"D3",x"E2",x"9A",x"86",x"01",x"4E",x"53",x"4B",x"B2",x"44",x"39",x"28",x"B6",x"1C",x"16",x"2F",x"6E",x"20",x"9D",x"66",x"B1",x"C6",x"9B",x"81",x"54",x"9A",x"65",x"EF",x"64",x"0A",x"96",x"75",x"56",x"2D",x"EA",x"28",x"84",x"CF",x"69",x"8E",x"4C",x"AC",x"30",x"91",x"B7",x"70",x"D2",x"B1",x"21",x"E4",x"28",x"25",x"AF",x"24",x"86",x"36",x"73",x"0A",x"C9",x"E2",x"18",x"56",x"DF",x"6B",x"52",x"51",x"6C",x"78",x"35",x"6F",x"54",x"D4",x"A6",x"12",x"65",x"DF",x"16",x"0E",x"4B",x"4A",x"96",x"75",x"C7",x"D8",x"62",x"2B",x"5D",x"D4",x"1B",x"65",x"4D",x"A5",x"1C",x"D1",x"37",x"99",x"BD",x"89",x"F2",x"59",x"BE",x"0C",x"35",x"D9",x"2A",x"11",x"63",x"5D",x"C8",x"9C",x"B0",x"9C",x"8D",x"4B",x"23",x"73",x"42",x"6A",x"63",x"67",x"5A",x"29",x"F1",x"03",x"FF",
		x"60",x"8C",x"32",x"79",x"CD",x"D8",x"DA",x"30",x"4C",x"D4",x"23",x"CB",x"6C",x"AA",x"10",x"B1",x"4A",x"AD",x"A2",x"8B",x"81",x"C5",x"2D",x"CB",x"CA",x"C4",x"0E",x"16",x"3B",x"B3",x"2A",x"6B",x"3A",x"58",x"DC",x"B4",x"8E",x"4C",x"EC",x"60",x"71",x"DC",x"D3",x"33",x"8E",x"43",x"CC",x"72",x"B5",x"88",x"AE",x"01",x"F5",x"AB",x"94",x"4D",x"5B",x"05",x"D4",x"F7",x"52",x"2A",x"69",x"E7",x"50",x"D3",x"4B",x"B8",x"BC",x"AB",x"41",x"6D",x"6F",x"A6",x"8E",x"2C",x"0A",x"73",x"DB",x"82",x"B8",x"66",x"1B",x"DC",x"CE",x"56",x"11",x"6D",x"6D",x"70",x"DB",x"CB",x"95",x"74",x"93",x"C1",x"75",x"A9",x"08",x"B4",x"D5",x"86",x"30",x"2D",x"DD",x"58",x"56",x"29",x"4A",x"D6",x"32",x"31",x"6F",x"C9",x"58",x"95",x"9A",x"39",x"22",x"0B",x"E3",x"58",x"EA",x"50",x"B5",x"2C",x"4A",x"32",x"B9",x"C2",x"59",x"5A",x"0B",x"D3",x"E4",x"31",x"F6",x"C8",x"A2",x"3C",x"E3",x"BA",x"CC",x"D9",x"33",x"0B",x"BD",x"ED",x"52",x"23",x"2F",x"22",x"72",x"B5",x"5D",x"58",x"B2",x"90",x"D8",x"A6",x"09",x"65",x"76",x"FB",x"00",x"FF",
		x"60",x"6D",x"2C",x"C2",x"A7",x"84",x"D7",x"AE",x"AE",x"72",x"ED",x"31",x"5C",x"B3",x"DA",x"CC",x"7D",x"5A",x"70",x"ED",x"6A",x"13",x"CF",x"19",x"85",x"25",x"AD",x"4B",x"24",x"67",x"12",x"96",x"84",x"BE",x"50",x"F6",x"75",x"88",x"E2",x"A6",x"CC",x"38",x"87",x"31",x"6A",x"58",x"0A",x"95",x"68",x"96",x"28",x"6E",x"2D",x"D8",x"A2",x"89",x"2A",x"AB",x"3D",x"C2",x"F0",x"11",x"8F",x"CA",x"AE",x"C0",x"DC",x"C2",x"D2",x"CE",x"03",x"FF",
		x"60",x"AE",x"4D",x"CE",x"C6",x"19",x"9C",x"84",x"39",x"B4",x"29",x"52",x"6C",x"93",x"76",x"EF",x"B3",x"C4",x"B0",x"4D",x"68",x"BC",x"CF",x"62",x"C7",x"76",x"69",x"F7",x"D1",x"53",x"05",x"DB",x"86",x"39",x"06",x"1D",x"17",x"48",x"E2",x"8E",x"10",x"A3",x"43",x"C1",x"B1",x"6A",x"43",x"EE",x"0A",x"03",x"26",x"A6",x"CE",x"16",x"A3",x"02",x"D4",x"86",x"32",x"5A",x"C9",x"08",x"68",x"E3",x"62",x"1F",x"35",x"4D",x"A1",x"8B",x"2B",x"63",x"34",x"F7",x"04",x"AF",x"6E",x"8D",x"5D",x"BD",x"0C",x"D8",x"85",x"CD",x"15",x"53",x"69",x"4A",x"E7",x"36",x"5F",x"5D",x"B8",x"45",x"59",x"58",x"7D",x"65",x"B1",x"21",x"67",x"61",x"8E",x"53",x"45",x"9B",x"A4",x"A9",x"3D",x"2D",x"63",x"D1",x"24",x"F2",x"00",x"FF",
		x"60",x"A6",x"AD",x"D2",x"DB",x"CC",x"E2",x"8C",x"BA",x"72",x"EF",x"0C",x"CA",x"B6",x"9A",x"2C",x"73",x"DC",x"A5",x"CB",x"AA",x"B3",x"CC",x"35",x"E3",x"AE",x"AB",x"8A",x"AE",x"DB",x"C4",x"D6",x"AC",x"2A",x"EA",x"EE",x"14",x"ED",x"BA",x"EA",x"CC",x"7B",x"D2",x"B0",x"EB",x"EA",x"2A",x"F3",x"9E",x"41",x"E7",x"63",x"28",x"DC",x"66",x"0A",x"D5",x"97",x"29",x"A8",x"DA",x"72",x"C8",x"1A",x"46",x"6F",x"7A",x"9C",x"29",x"B3",x"99",x"65",x"DA",x"72",x"D4",x"56",x"62",x"D1",x"B6",x"3B",x"58",x"52",x"3F",x"FF",
		x"60",x"21",x"88",x"22",x"27",x"14",x"BD",x"B6",x"30",x"B2",x"E8",x"76",x"E4",x"D6",x"92",x"60",x"7C",x"93",x"B1",x"75",x"49",x"6D",x"C8",x"35",x"B4",x"4E",x"29",x"93",x"AD",x"0B",x"C5",x"3B",x"B5",x"DC",x"EB",x"D8",x"50",x"E8",x"5C",x"2A",x"AF",x"62",x"D3",x"C0",x"4F",x"6A",x"23",x"F7",x"0D",x"03",x"2D",x"A6",x"D7",x"BA",x"97",x"59",x"3C",x"99",x"81",x"87",x"E9",x"60",x"71",x"AD",x"66",x"5A",x"66",x"92",x"25",x"35",x"59",x"58",x"DA",x"0C",x"51",x"39",x"0F",x"FF",
		x"60",x"21",x"8B",x"2E",x"CA",x"85",x"33",x"37",x"2F",x"B8",x"0A",x"33",x"EE",x"5A",x"6C",x"1B",x"C3",x"D5",x"64",x"73",x"72",x"4C",x"0C",x"33",x"B6",x"AE",x"C9",x"F6",x"C3",x"84",x"DD",x"5A",x"27",x"C7",x"77",x"13",x"65",x"EB",x"92",x"3C",x"5F",x"34",x"0D",x"B9",x"4B",x"F2",x"6D",x"0D",x"63",x"E7",x"2E",x"29",x"54",x"DE",x"33",x"92",x"D2",x"85",x"48",x"EB",x"4C",x"6B",x"49",x"EA",x"72",x"97",x"2D",x"4C",x"29",x"AD",x"AB",x"9D",x"F7",x"08",x"47",x"6F",x"6C",x"D4",x"35",x"D4",x"44",x"B2",x"3E",x"FF",
		x"60",x"C5",x"C8",x"3C",x"47",x"C5",x"16",x"17",x"2F",x"E9",x"6A",x"52",x"BF",x"34",x"D2",x"C2",x"A3",x"D5",x"AC",x"76",x"CB",x"92",x"EB",x"62",x"F6",x"D9",x"A5",x"48",x"BE",x"9B",x"45",x"6B",x"97",x"2A",x"A4",x"0C",x"AC",x"2E",x"33",x"EA",x"2C",x"63",x"44",x"ED",x"C9",x"A8",x"32",x"F7",x"75",x"97",x"D7",x"A3",x"CB",x"DC",x"47",x"4C",x"5F",x"8F",x"A1",x"73",x"99",x"70",x"DA",x"32",x"C6",x"4A",x"65",x"33",x"79",x"4B",x"9B",x"82",x"AE",x"E1",x"88",x"C7",x"6D",x"09",x"AE",x"8A",x"22",x"2F",x"A7",x"35",x"F8",x"6A",x"F2",x"BA",x"18",x"B6",x"60",x"B3",x"31",x"6A",x"94",x"D8",x"A2",x"8E",x"61",x"A9",x"39",x"0F",x"FF",
		x"60",x"8E",x"49",x"26",x"32",x"38",x"6A",x"15",x"39",x"F8",x"48",x"B5",x"B8",x"53",x"8C",x"A0",x"B2",x"D4",x"F5",x"56",x"B2",x"7D",x"0C",x"E5",x"C9",x"D1",x"C5",x"0E",x"CE",x"5D",x"CC",x"9F",x"34",x"3B",x"B8",x"70",x"76",x"7B",x"92",x"2C",x"15",x"A3",x"CC",x"F3",x"52",x"B2",x"64",x"9C",x"94",x"F1",x"D9",x"C1",x"12",x"69",x"CA",x"D3",x"2E",x"07",x"5B",x"D9",x"E9",x"4C",x"BA",x"9D",x"1C",x"63",x"27",x"68",x"63",x"76",x"70",x"9D",x"9A",x"A4",x"F1",x"29",x"CE",x"B5",x"AA",x"CA",x"8B",x"2F",x"07",x"D7",x"E9",x"2A",x"2E",x"9B",x"1C",x"5C",x"AF",x"AA",x"2D",x"65",x"76",x"70",x"83",x"4B",x"A7",x"B0",x"DB",x"C1",x"0D",x"3E",x"9D",x"C2",x"2F",x"27",x"2F",x"71",x"6F",x"0B",x"5C",x"1C",x"BC",x"68",x"3A",x"A0",x"63",x"72",x"F0",x"83",x"EC",x"A6",x"F2",x"49",x"C1",x"CF",x"4C",x"BB",x"16",x"EA",x"84",x"C0",x"9B",x"2A",x"4D",x"BB",x"98",x"42",x"EB",x"3B",x"B9",x"E3",x"76",x"8A",x"82",x"CC",x"F6",x"94",x"27",x"29",x"0A",x"2A",x"DA",x"53",x"1E",x"97",x"38",x"AB",x"48",x"71",x"79",x"93",x"D2",x"AC",x"A2",x"D4",x"68",x"49",x"4A",x"92",x"CB",x"64",x"95",x"25",x"21",x"C9",x"36",x"52",x"94",x"9E",x"86",x"34",x"D9",x"48",x"51",x"99",x"E3",x"B2",x"50",x"4D",x"25",x"AB",x"B2",x"CB",x"42",x"71",x"A5",x"AC",x"09",x"2E",x"0F",x"CD",x"44",x"AA",x"4B",x"BA",x"C2",x"E4",x"0C",x"8B",x"98",x"68",x"0A",x"53",x"C3",x"AD",x"6A",x"A4",x"29",x"74",x"A9",x"D0",x"CC",x"89",x"A6",x"72",x"21",x"53",x"3D",x"6E",x"9A",x"3A",x"6A",x"4F",x"51",x"5B",x"C4",x"BA",x"A0",x"A2",x"42",x"2D",x"E1",x"03",x"FF",
		x"60",x"6D",x"9F",x"96",x"3D",x"5B",x"D4",x"B6",x"25",x"D9",x"28",x"15",x"D9",x"B2",x"D6",x"A6",x"39",x"CB",x"D9",x"EB",x"3A",x"A2",x"F2",x"76",x"93",x"3D",x"AB",x"AF",x"42",x"AA",x"92",x"B3",x"9E",x"A5",x"0B",x"89",x"0E",x"F1",x"77",x"E6",x"61",x"C4",x"AB",x"98",x"5B",x"E9",x"8B",x"F2",x"0A",x"A1",x"7E",x"A1",x"8F",x"26",x"DA",x"C4",x"F7",x"B4",x"A5",x"71",x"A9",x"4C",x"F5",x"32",x"C6",x"61",x"D5",x"26",x"99",x"EB",x"98",x"1B",x"57",x"DF",x"30",x"3D",x"E7",x"18",x"52",x"22",x"8B",x"DD",x"8D",x"BD",x"4B",x"F6",x"6E",x"D5",x"BA",x"D6",x"2E",x"38",x"A6",x"C5",x"DD",x"98",x"BB",x"C6",x"EC",x"73",x"67",x"6B",x"5F",x"56",x"AD",x"53",x"99",x"AD",x"6D",x"1B",x"95",x"AA",x"40",x"5F",x"8E",x"2E",x"39",x"AB",x"D8",x"4B",x"D8",x"23",x"9F",x"3A",x"D7",x"2C",x"0F",x"FF",
		x"60",x"C1",x"0E",x"2D",x"D5",x"7C",x"4A",x"17",x"35",x"C6",x"76",x"93",x"1A",x"D5",x"E4",x"68",x"D7",x"24",x"7C",x"72",x"93",x"83",x"1F",x"33",x"8B",x"59",x"4D",x"09",x"6E",x"5C",x"CD",x"67",x"37",x"3D",x"E8",x"CE",x"10",x"79",x"54",x"6C",x"EF",x"C6",x"8C",x"7D",x"96",x"F3",x"7C",x"19",x"55",x"CE",x"D3",x"26",x"50",x"65",x"D5",x"35",x"47",x"AB",x"48",x"AD",x"64",x"CF",x"AE",x"CD",x"62",x"51",x"C7",x"D4",x"32",x"D6",x"03",x"FF",
		x"60",x"4C",x"16",x"BD",x"45",x"23",x"6C",x"35",x"AD",x"63",x"89",x"0E",x"8E",x"DD",x"3C",x"AF",x"27",x"D1",x"73",x"65",x"B2",x"83",x"EC",x"86",x"CC",x"56",x"41",x"0D",x"6A",x"0A",x"32",x"1B",x"1A",x"CE",x"F1",x"1A",x"74",x"EB",x"22",x"68",x"52",x"AE",x"D5",x"2D",x"35",x"23",x"58",x"DE",x"30",x"37",x"27",x"0F",x"FF",
		x"60",x"C6",x"69",x"4C",x"C4",x"BA",x"4B",x"36",x"BB",x"3B",x"43",x"89",x"A9",x"D3",x"CC",x"AE",x"0C",x"35",x"7B",x"E2",x"30",x"BA",x"73",x"94",x"AE",x"9A",x"43",x"6F",x"52",x"D0",x"BB",x"22",x"0F",x"A3",x"5B",x"43",x"89",x"A9",x"CD",x"6C",x"2F",x"C4",x"76",x"CA",x"32",x"30",x"20",x"51",x"CB",x"14",x"0F",x"23",x"C2",x"DE",x"8D",x"4A",x"54",x"B5",x"30",x"47",x"37",x"6A",x"71",x"89",x"C4",x"99",x"D9",x"69",x"C4",x"31",x"88",x"56",x"44",x"D7",x"91",x"C5",x"64",x"52",x"2E",x"9D",x"5B",x"EE",x"AB",x"4B",x"A7",x"6E",x"2E",x"4D",x"AC",x"C1",x"15",x"D2",x"19",x"45",x"B5",x"86",x"9B",x"AA",x"65",x"96",x"54",x"E3",x"EE",x"EA",x"4E",x"59",x"5A",x"94",x"9B",x"7B",x"38",x"45",x"40",x"74",x"11",x"04",x"C8",x"2E",x"9D",x"01",x"C9",x"A9",x"A7",x"2A",x"69",x"B7",x"B0",x"70",x"DC",x"CA",x"E8",x"B4",x"54",x"B5",x"CB",x"A8",x"92",x"55",x"4F",x"D6",x"BE",x"A3",x"8E",x"C6",x"C2",x"4C",x"F3",x"8E",x"26",x"59",x"0D",x"55",x"C9",x"33",x"BA",x"64",x"23",x"44",x"44",x"6F",x"EB",x"93",x"B2",x"70",x"53",x"7D",x"6D",x"C8",x"C6",x"C2",x"9D",x"F4",x"95",x"31",x"1B",x"4F",x"35",x"D4",x"56",x"A6",x"AC",x"D5",x"35",x"D9",x"2F",x"9A",x"92",x"17",x"53",x"37",x"AF",x"6E",x"8E",x"56",x"C2",x"4D",x"33",x"9B",x"36",x"59",x"0F",x"51",x"F6",x"67",x"FA",x"AC",x"CC",x"C3",x"44",x"1F",x"20",x"80",x"47",x"CF",x"12",x"15",x"2B",x"A6",x"9E",x"B5",x"5B",x"58",x"92",x"18",x"7B",x"B7",x"6E",x"41",x"0C",x"16",x"61",x"3D",x"BB",x"F9",x"D1",x"56",x"98",x"D9",x"A3",x"E6",x"45",x"D3",x"A5",x"AA",x"AD",x"8A",x"EB",x"4D",x"37",x"BB",x"C6",x"4E",x"AE",x"B5",x"31",x"AC",x"EE",x"38",x"F8",x"41",x"45",x"3A",x"51",x"5D",x"14",x"E7",x"C0",x"C6",x"5E",x"8D",x"18",x"50",x"4C",x"AA",x"00",x"9A",x"36",x"63",x"C0",x"CC",x"A6",x"0C",x"98",x"77",x"5C",x"00",x"63",x"47",x"28",x"60",x"CC",x"4A",x"01",x"8C",x"91",x"29",x"80",x"3E",x"23",x"4A",x"51",x"23",x"89",x"64",x"B6",x"19",x"65",x"71",x"6C",x"EA",x"D6",x"6D",x"34",x"55",x"AB",x"B9",x"8B",x"FB",x"D1",x"15",x"A5",x"11",x"4E",x"CE",x"47",x"57",x"8C",x"B8",x"A6",x"38",x"17",x"40",x"8B",x"16",x"A3",x"E9",x"D1",x"0C",x"55",x"96",x"8D",x"AA",x"5B",x"35",x"F6",x"58",x"D5",x"B2",x"AA",x"55",x"5D",x"67",x"55",x"08",x"8A",x"11",x"53",x"BF",x"58",x"04",x"90",x"21",x"82",x"00",x"D6",x"B9",x"21",x"20",x"1A",x"93",x"07",x"FF",
		x"60",x"42",x"4E",x"54",x"2D",x"BB",x"A3",x"24",x"A9",x"31",x"A5",x"E8",x"28",x"5C",x"A4",x"1A",x"58",x"52",x"7D",x"64",x"93",x"8A",x"35",x"0D",x"E3",x"4B",x"45",x"8E",x"29",x"58",x"5C",x"27",x"25",x"2D",x"64",x"35",x"65",x"5F",x"E4",x"9C",x"14",x"30",x"54",x"D2",x"89",x"C9",x"B3",x"10",x"8E",x"CA",x"2A",x"04",x"98",x"89",x"4D",x"00",x"6B",x"A6",x"09",x"60",x"0E",x"E7",x"11",x"17",x"A7",x"6C",x"91",x"4B",x"46",x"92",x"6D",x"48",x"64",x"AC",x"1E",x"79",x"D6",x"A3",x"9E",x"B1",x"68",x"D4",x"D9",x"B4",x"B9",x"E5",x"E5",x"D2",x"15",x"5D",x"E6",x"96",x"77",x"18",x"50",x"AC",x"39",x"03",x"AA",x"51",x"65",x"40",x"36",x"C1",x"26",x"6B",x"22",x"C3",x"3C",x"96",x"B8",x"6A",x"28",x"CB",x"08",x"DD",x"EC",x"BA",x"21",x"22",x"CD",x"BC",x"AD",x"00",x"86",x"66",x"55",x"C0",x"4A",x"29",x"02",x"98",x"3B",x"2D",x"65",x"D9",x"93",x"65",x"66",x"ED",x"56",x"E5",x"A0",x"11",x"1E",x"4B",x"5A",x"97",x"63",x"94",x"AB",x"2F",x"69",x"6D",x"8E",x"D5",x"9C",x"31",x"A7",x"D5",x"39",x"D4",x"A8",x"C6",x"92",x"54",x"E5",x"D0",x"E9",x"1A",x"77",x"08",x"E0",x"9B",x"19",x"02",x"7C",x"D6",x"00",x"04",x"84",x"1E",x"41",x"80",x"D8",x"23",x"87",x"93",x"5C",x"88",x"6B",x"57",x"1E",x"4E",x"72",x"5A",x"2E",x"5D",x"25",x"B9",x"21",x"B9",x"9B",x"64",x"55",x"00",x"60",x"40",x"71",x"69",x"04",x"90",x"29",x"22",x"19",x"3E",x"76",x"A8",x"68",x"99",x"A2",x"85",x"1E",x"CE",x"3E",x"41",x"8B",x"1A",x"C2",x"86",x"A8",x"8D",x"29",x"4A",x"28",x"6D",x"A2",x"3E",x"B5",x"28",x"3E",x"A7",x"8B",x"D5",x"D4",x"22",x"7A",x"1F",x"69",x"12",x"8B",x"92",x"9C",x"1C",x"95",x"6A",x"D4",x"54",x"40",x"2B",x"EA",x"0A",x"68",x"C9",x"CC",x"A8",x"CD",x"49",x"56",x"B8",x"14",x"A3",x"54",x"A3",x"16",x"11",x"B1",x"4B",x"5A",x"23",x"99",x"79",x"34",x"69",x"79",x"8A",x"6C",x"96",x"B9",x"78",x"94",x"D5",x"A4",x"51",x"46",x"D3",x"D1",x"0F",x"E5",x"49",x"A6",x"6B",x"C3",x"5C",x"85",x"A8",x"BB",x"D6",x"71",x"73",x"55",x"A4",x"A1",x"5E",x"C7",x"AD",x"CD",x"A0",x"B9",x"79",x"5C",x"B7",x"25",x"2B",x"A6",x"D1",x"4D",x"C2",x"5A",x"4C",x"28",x"55",x"36",x"79",x"FF",
		x"60",x"A6",x"AE",x"82",x"55",x"3A",x"1B",x"B9",x"26",x"5A",x"92",x"DE",x"48",x"94",x"AA",x"10",x"C9",x"DD",x"63",x"75",x"AB",x"A2",x"4E",x"8B",x"90",x"6C",x"AD",x"8A",x"BA",x"DD",x"0A",x"BB",x"B6",x"2A",x"B8",x"D6",x"6C",x"E8",x"5C",x"AA",x"10",x"4B",x"A2",x"61",x"73",x"A9",x"63",x"73",x"CA",x"A2",x"5C",x"A9",x"CC",x"1B",x"A5",x"55",x"3B",x"32",x"A0",x"8E",x"30",x"06",x"8C",x"51",x"C6",x"80",x"D9",x"D3",x"19",x"30",x"73",x"1A",x"03",x"46",x"AF",x"68",x"51",x"6F",x"26",x"A6",x"92",x"74",x"A4",x"29",x"5B",x"9A",x"F5",x"DC",x"91",x"67",x"5D",x"55",x"26",x"73",x"47",x"99",x"4D",x"57",x"98",x"3C",x"1D",x"75",x"B6",x"5D",x"E1",x"B2",x"64",x"D4",x"C5",x"4D",x"B8",x"F9",x"9D",x"D1",x"66",x"5B",x"1A",x"32",x"73",x"41",x"00",x"39",x"44",x"31",x"20",x"EB",x"2A",x"06",x"54",x"55",x"C9",x"80",x"26",x"A6",x"08",x"10",x"45",x"05",x"CB",x"3D",x"8B",x"C8",x"74",x"DB",x"AA",x"D2",x"CA",x"33",x"35",x"23",x"B7",x"B2",x"06",x"75",x"B2",x"AE",x"32",x"F2",x"9A",x"3C",x"D4",x"72",x"CE",x"C8",x"4B",x"C9",x"30",x"CF",x"2A",x"23",x"2F",x"BE",x"22",x"3C",x"E6",x"8C",x"2C",x"FB",x"AA",x"94",x"98",x"D3",x"B2",x"98",x"DB",x"CD",x"6B",x"4A",x"CB",x"62",x"1E",x"17",x"AD",x"C9",x"2D",x"F3",x"A9",x"42",x"2D",x"E3",x"B6",x"34",x"7A",x"2B",x"D1",x"88",x"5A",x"F2",x"6A",x"DB",x"35",x"AC",x"B4",x"00",x"8A",x"E8",x"64",x"40",x"16",x"1B",x"0C",x"48",x"66",x"82",x"01",x"49",x"75",x"12",x"20",x"91",x"69",x"04",x"C8",x"AE",x"0E",x"02",x"C8",x"DC",x"AD",x"79",x"C9",x"BB",x"59",x"66",x"95",x"16",x"86",x"E6",x"1A",x"5D",x"65",x"5B",x"1C",x"F3",x"28",x"67",x"55",x"69",x"69",x"F6",x"E7",x"14",x"51",x"A7",x"E5",x"C5",x"AC",x"B3",x"C7",x"EC",x"56",x"15",x"B3",x"C6",x"11",x"93",x"5B",x"5D",x"6D",x"B9",x"48",x"4C",x"6E",x"75",x"32",x"1A",x"66",x"15",x"BB",x"94",x"D1",x"87",x"AB",x"A5",x"E9",x"52",x"26",x"97",x"26",x"EA",x"61",x"46",x"5D",x"6D",x"86",x"B1",x"97",x"19",x"5D",x"09",x"E9",x"1A",x"31",x"7B",x"34",x"25",x"78",x"6A",x"46",x"ED",x"91",x"66",x"9F",x"61",x"DE",x"B5",x"47",x"5C",x"6C",x"84",x"CB",x"CC",x"09",x"59",x"D5",x"A9",x"86",x"56",x"99",x"01",x"CA",x"85",x"95",x"30",x"B8",x"E4",x"A8",x"9C",x"9D",x"C2",x"50",x"28",x"2A",x"73",x"51",x"8A",x"42",x"21",x"CF",x"F0",x"26",x"31",x"72",x"A1",x"CB",x"62",x"11",x"6E",x"07",x"80",x"00",x"C9",x"58",x"BA",x"38",x"78",x"57",x"9D",x"8A",x"D3",x"A2",x"10",x"C6",x"C5",x"6A",x"CA",x"48",x"A2",x"6B",x"33",x"AB",x"C9",x"23",x"CD",x"C9",x"4D",x"35",x"67",x"8F",x"AC",x"44",x"55",x"8B",x"5C",x"3C",x"8A",x"5A",x"54",x"34",x"B2",x"F5",x"A8",x"6B",x"51",x"E6",x"F2",x"2D",x"A3",x"A9",x"C5",x"98",x"D3",x"B6",x"8C",x"B2",x"64",x"96",x"28",x"6F",x"D3",x"A6",x"32",x"44",x"C2",x"65",x"49",x"9B",x"72",x"17",x"89",x"92",x"B5",x"65",x"C9",x"83",x"D5",x"DD",x"9A",x"A5",x"2D",x"0F",x"31",x"35",x"6D",x"97",x"F6",x"D2",x"4C",x"D5",x"79",x"69",x"3A",x"4B",x"52",x"D1",x"90",x"2E",x"E6",x"C8",x"45",x"44",x"43",x"DB",x"22",x"40",x"67",x"6A",x"02",x"84",x"68",x"42",x"80",x"A4",x"8B",x"11",x"10",x"6D",x"08",x"02",x"92",x"48",x"45",x"40",x"E4",x"2D",x"0F",x"FF",
		x"60",x"08",x"C8",x"CE",x"95",x"00",x"35",x"84",x"12",x"20",x"1B",x"F3",x"12",x"C5",x"41",x"19",x"A6",x"4D",x"5A",x"98",x"06",x"7B",x"BA",x"74",x"69",x"51",x"9E",x"9C",x"AE",x"B1",x"6A",x"84",x"A5",x"A8",x"59",x"E4",x"EC",x"11",x"D6",x"E8",x"EA",x"D6",x"75",x"46",x"54",x"9C",x"8B",x"C7",x"54",x"19",x"71",x"D1",x"85",x"E1",x"55",x"B5",x"A5",x"D9",x"9A",x"B8",x"AC",x"E2",x"96",x"A7",x"A8",x"CE",x"56",x"AA",x"5B",x"95",x"0A",x"AB",x"4B",x"BA",x"6A",x"75",x"4E",x"AC",x"6A",x"19",x"A9",x"35",x"C5",x"99",x"B8",x"55",x"68",x"03",x"34",x"DD",x"22",x"80",x"92",x"16",x"41",x"00",x"D1",x"AA",x"B7",x"B2",x"45",x"0C",x"B1",x"8D",x"35",x"EA",x"12",x"54",x"39",x"6A",x"76",x"E9",x"92",x"A4",x"2C",x"49",x"5B",x"A9",x"4B",x"82",x"62",x"2C",x"22",x"A7",x"2E",x"4A",x"2A",x"97",x"8A",x"1C",x"FA",x"A2",x"31",x"CC",x"D3",x"B6",x"00",x"9A",x"66",x"55",x"C0",x"68",x"93",x"AD",x"C9",x"99",x"4C",x"BD",x"92",x"B6",x"2A",x"16",x"4E",x"B5",x"5A",x"32",x"EA",x"68",x"2B",x"C2",x"69",x"D3",x"A8",x"82",x"D9",x"52",x"D5",x"D6",x"A3",x"8C",x"E6",x"8A",x"D5",x"53",x"8F",x"3C",x"FA",x"49",x"15",x"5F",x"34",x"B2",x"58",x"DA",x"44",x"A3",x"D6",x"48",x"62",x"31",x"B3",x"CC",x"DA",x"23",x"AE",x"91",x"43",x"3C",x"66",x"B7",x"B8",x"65",x"56",x"89",x"AA",x"55",x"92",x"64",x"24",x"CB",x"CD",x"4C",x"49",x"A2",x"C9",x"08",x"E1",x"D8",x"23",x"6E",x"4E",x"39",x"A3",x"82",x"8C",x"A8",x"5A",x"E5",x"8A",x"08",x"37",x"C2",x"62",x"45",x"32",x"2B",x"EC",x"08",x"8B",x"63",x"F5",x"EA",x"28",x"23",x"28",x"9E",x"5D",x"7B",x"6C",x"B5",x"20",x"59",x"95",x"CC",x"36",x"1D",x"7C",x"AF",x"B5",x"34",x"4B",x"76",x"F2",x"A2",x"16",x"4F",x"2F",x"2B",x"C9",x"8B",x"9A",x"23",x"A2",x"A4",x"24",x"2F",x"1A",x"8E",x"CC",x"94",x"52",x"FC",x"EC",x"59",x"22",x"D3",x"4C",x"0A",x"92",x"56",x"F7",x"2A",x"29",x"2E",x"CC",x"4E",x"D4",x"AB",x"A5",x"08",x"3F",x"29",x"71",x"8B",x"96",x"22",x"BC",x"64",x"C4",x"3C",x"8B",x"0E",x"F3",x"82",x"34",x"8F",x"28",x"D3",x"CC",x"F3",x"DA",x"2D",x"32",x"2C",x"B7",x"A4",x"55",x"33",x"C9",x"8A",x"33",x"E2",x"56",x"54",x"25",x"26",x"CE",x"08",x"5A",x"10",x"E3",x"1A",x"DB",x"C1",x"F7",x"C6",x"B2",x"B8",x"99",x"8C",x"A0",x"19",x"D2",x"88",x"0A",x"3D",x"92",x"6E",x"99",x"AD",x"27",x"F4",x"C8",x"BB",x"50",x"F4",x"E9",x"52",x"A3",x"1E",x"CA",x"40",x"B2",x"66",x"B7",x"AE",x"39",x"01",x"F3",x"2E",x"63",x"FA",x"6E",x"4D",x"CC",x"26",x"96",x"00",x"AE",x"52",x"11",x"C0",x"0C",x"A9",x"65",x"E8",x"C6",x"C5",x"2C",x"6A",x"97",x"21",x"5B",x"B3",x"B4",x"2C",x"DD",x"86",x"E8",x"CA",x"C3",x"AA",x"72",x"1B",x"63",x"2A",x"0D",x"CF",x"B2",x"63",x"8A",x"B9",x"C4",x"33",x"CA",x"B4",x"29",x"D9",x"13",x"3E",x"B7",x"3C",x"E6",x"98",x"CB",x"DC",x"B3",x"CC",x"58",x"72",x"0A",x"37",x"EB",x"B2",x"63",x"CB",x"D5",x"5D",x"63",x"A2",x"8E",x"BD",x"86",x"36",x"F7",x"1C",x"3B",x"8E",x"9A",x"DD",x"35",x"B2",x"72",x"3B",x"6A",x"51",x"97",x"AC",x"C8",x"6D",x"6A",x"D9",x"54",x"AD",x"A2",x"94",x"B1",x"46",x"17",x"8F",x"08",x"5B",x"A6",x"9A",x"C3",x"54",x"B3",x"4A",x"98",x"73",x"F2",x"50",x"AD",x"D0",x"E1",x"2C",x"21",x"CD",x"C4",x"CB",x"3C",x"FF",
		x"60",x"62",x"B0",x"3C",x"B2",x"CC",x"AC",x"98",x"4E",x"6A",x"6F",x"17",x"B7",x"5D",x"B2",x"AC",x"A4",x"2C",x"D3",x"F2",x"08",x"4B",x"16",x"B7",x"2E",x"C7",x"C3",x"2D",x"DD",x"5D",x"B3",x"AC",x"0C",x"2B",x"37",x"0B",x"CD",x"B2",x"DB",x"F4",x"DC",x"DC",x"BC",x"22",x"5A",x"53",x"D2",x"74",x"B3",x"8E",x"30",x"4D",x"49",x"2D",x"4D",x"C7",x"83",x"35",x"3D",x"D6",x"32",x"ED",x"A8",x"D2",x"DC",x"D8",x"C2",x"AC",x"A2",x"6A",x"0B",x"42",x"37",x"F7",x"8C",x"78",x"A5",x"09",x"31",x"CA",x"2C",x"A3",x"84",x"21",x"56",x"B7",x"6C",x"B7",x"22",x"80",x"D4",x"42",x"CB",x"98",x"AB",x"B9",x"67",x"84",x"6D",x"53",x"AE",x"12",x"5D",x"6A",x"77",x"0C",x"39",x"4B",x"44",x"79",x"D4",x"31",x"E6",x"C2",x"E9",x"DD",x"51",x"C6",x"54",x"7C",x"AA",x"77",x"CE",x"19",x"53",x"75",x"A5",x"56",x"39",x"67",x"CC",x"C5",x"97",x"5A",x"E5",x"9C",x"31",x"15",x"57",x"66",x"19",x"73",x"C6",x"54",x"6C",x"9B",x"56",x"CC",x"19",x"63",x"31",x"6D",x"96",x"31",x"7B",x"F4",x"C5",x"94",x"B9",x"E5",x"9D",x"D6",x"65",x"9B",x"EA",x"D6",x"93",x"4B",x"1E",x"6C",x"6A",x"C5",x"96",x"49",x"91",x"F7",x"29",x"53",x"1D",x"3A",x"04",x"89",x"87",x"A6",x"F6",x"28",x"E7",x"27",x"9E",x"E2",x"5A",x"B3",x"19",x"90",x"54",x"1A",x"03",x"B2",x"4D",x"65",x"40",x"D1",x"A5",x"04",x"88",x"7C",x"0C",x"01",x"49",x"A6",x"3E",x"FF",
		x"60",x"AA",x"D7",x"71",x"D8",x"A2",x"62",x"9B",x"C6",x"96",x"C0",x"A8",x"B2",x"9D",x"F2",x"68",x"9A",x"D5",x"3B",x"CE",x"08",x"53",x"08",x"B1",x"98",x"A8",x"23",x"C8",x"2E",x"C4",x"A2",x"26",x"07",x"CF",x"5B",x"49",x"E7",x"AA",x"5D",x"DC",x"E8",x"C5",x"C4",x"A2",x"CE",x"F0",x"8A",x"33",x"35",x"EF",x"22",x"CE",x"4B",x"C6",x"34",x"6A",x"4C",x"03",x"03",x"9A",x"2C",x"2D",x"6E",x"65",x"A1",x"AE",x"59",x"B9",x"B9",x"C5",x"88",x"49",x"6D",x"D8",x"E6",x"15",x"2D",x"66",x"B1",x"65",x"86",x"57",x"A4",x"AA",x"FB",x"94",x"56",x"7E",x"D0",x"26",x"51",x"6D",x"18",x"85",x"56",x"86",x"67",x"97",x"A8",x"90",x"36",x"9D",x"A6",x"6A",x"56",x"4C",x"90",x"0D",x"A9",x"CF",x"59",x"75",x"6E",x"36",x"62",x"5A",x"1B",x"35",x"78",x"59",x"8B",x"59",x"6E",x"99",x"56",x"35",x"A3",x"EC",x"D1",x"95",x"47",x"D1",x"75",x"90",x"66",x"8D",x"0A",x"55",x"14",x"14",x"E5",x"59",x"26",x"34",x"51",x"60",x"57",x"A8",x"95",x"D6",x"B4",x"28",x"4E",x"A6",x"4D",x"4C",x"9E",x"B5",x"88",x"98",x"A6",x"15",x"79",x"D6",x"22",x"E6",x"9A",x"66",x"E4",x"25",x"99",x"B2",x"7B",x"E3",x"91",x"16",x"2B",x"A6",x"51",x"AB",x"47",x"5C",x"AC",x"9A",x"DA",x"CE",x"6E",x"61",x"D5",x"21",x"C6",x"55",x"A6",x"84",x"4B",x"85",x"A8",x"48",x"E2",x"E6",x"56",x"59",x"AC",x"56",x"95",x"86",x"93",x"BC",x"89",x"E5",x"94",x"29",x"5E",x"CA",x"AC",x"1A",x"39",x"05",x"25",x"C5",x"8A",x"A9",x"E7",x"A2",x"E6",x"E5",x"A0",x"A6",x"9A",x"4D",x"86",x"97",x"BC",x"B9",x"79",x"8E",x"19",x"5E",x"34",x"19",x"A6",x"5D",x"A5",x"F9",x"3E",x"B5",x"98",x"4F",x"94",x"12",x"46",x"93",x"EA",x"1E",x"66",x"53",x"6A",x"E3",x"70",x"86",x"5B",x"6B",x"85",x"F7",x"1D",x"22",x"53",x"BB",x"74",x"59",x"46",x"19",x"D5",x"62",x"04",x"44",x"67",x"5E",x"FA",x"AC",x"3D",x"55",x"2B",x"EE",x"18",x"BA",x"71",x"31",x"A9",x"D9",x"AD",x"AF",x"5E",x"59",x"72",x"EB",x"B4",x"A9",x"1B",x"15",x"F6",x"A9",x"55",x"96",x"A6",x"C5",x"AC",x"4B",x"4A",x"59",x"AB",x"34",x"B7",x"52",x"E5",x"61",x"EF",x"46",x"94",x"D3",x"A3",x"3E",x"FF",
		x"60",x"2B",x"EE",x"C1",x"43",x"22",x"96",x"AC",x"A0",x"86",x"54",x"CD",x"9C",x"BB",x"DC",x"9A",x"4C",x"D2",x"6B",x"76",x"72",x"6A",x"C3",x"70",x"EB",x"2A",x"04",x"48",x"9E",x"4C",x"00",x"B9",x"93",x"1B",x"A0",x"DB",x"73",x"05",x"4C",x"95",x"6A",x"82",x"16",x"D2",x"34",x"72",x"AE",x"F2",x"6A",x"74",x"C9",x"C8",x"2A",x"02",x"68",x"39",x"2D",x"39",x"B1",x"A0",x"57",x"E8",x"EA",x"66",x"85",x"2C",x"56",x"29",x"AB",x"9A",x"15",x"BB",x"69",x"B8",x"2F",x"6C",x"6E",x"2C",x"E9",x"E1",x"3E",x"2B",x"04",x"B1",x"47",x"98",x"E7",x"1C",x"28",x"75",x"18",x"15",x"16",x"3E",x"BB",x"C5",x"B1",x"76",x"B8",x"EB",x"AA",x"16",x"86",x"E9",x"11",x"16",x"0B",x"5B",x"10",x"47",x"6A",x"94",x"B5",x"6A",x"7E",x"1A",x"6E",x"99",x"BA",x"AA",x"05",x"B9",x"AB",x"57",x"C8",x"CA",x"16",x"E6",x"41",x"51",x"AE",x"8B",x"5C",x"1C",x"2A",x"56",x"8A",x"24",x"49",x"69",x"AC",x"AA",x"E1",x"6C",x"A5",x"64",x"A1",x"A9",x"A5",x"AB",x"ED",x"52",x"A7",x"C9",x"56",x"C9",x"A9",x"CA",x"90",x"06",x"6B",x"0E",x"A7",x"2A",x"53",x"5A",x"AC",x"59",x"DC",x"2A",x"AD",x"F9",x"90",x"A7",x"EB",x"A2",x"B0",x"A6",x"83",x"DE",x"49",x"BD",x"DD",x"96",x"0E",x"44",x"07",x"6F",x"76",x"7B",x"BA",x"10",x"ED",x"D2",x"D9",x"1D",x"F9",x"90",x"57",x"48",x"16",x"75",x"A6",x"21",x"9C",x"6D",x"6E",x"1E",x"FF",
		x"60",x"6D",x"2F",x"46",x"D3",x"BA",x"6A",x"8F",x"B1",x"47",x"4B",x"71",x"5F",x"3A",x"FA",x"9A",x"3D",x"39",x"F4",x"69",x"1B",x"5A",x"D3",x"90",x"90",x"25",x"04",x"08",x"91",x"9A",x"01",x"A5",x"95",x"0A",x"20",x"25",x"57",x"03",x"0C",x"19",x"9A",x"DA",x"65",x"2B",x"D4",x"24",x"6B",x"E8",x"5B",x"F2",x"64",x"B7",x"35",x"A6",x"6F",x"CD",x"92",x"43",x"56",x"33",x"20",x"44",x"D6",x"52",x"A7",x"4C",x"6E",x"21",x"AB",x"47",x"55",x"2A",x"99",x"9B",x"76",x"19",x"65",x"09",x"21",x"6E",x"B6",x"76",x"E4",x"39",x"84",x"B8",x"F7",x"9C",x"51",x"54",x"15",x"E2",x"96",x"93",x"15",x"30",x"89",x"A9",x"00",x"96",x"2C",x"17",x"C0",x"C2",x"E2",x"02",x"38",x"3A",x"4A",x"01",x"25",x"B9",x"80",x"00",x"4A",x"50",x"19",x"41",x"1B",x"2E",x"CA",x"9C",x"7A",x"04",x"2D",x"19",x"B2",x"D7",x"EA",x"E1",x"0D",x"EB",x"4C",x"56",x"AB",x"87",x"3B",x"42",x"12",x"6A",x"35",x"1E",x"EE",x"B4",x"C1",x"A8",x"D5",x"66",x"F8",x"D3",x"17",x"13",x"E7",x"92",x"11",x"4E",x"17",x"44",x"5A",x"4B",x"46",x"34",x"42",x"20",x"79",x"CD",x"19",x"49",x"8B",x"02",x"9A",x"53",x"77",x"64",x"5D",x"29",x"6A",x"76",x"A3",x"91",x"37",x"A9",x"A8",x"33",x"B5",x"47",x"D5",x"83",x"21",x"6B",x"2F",x"19",x"4D",x"8F",x"01",x"A4",x"B5",x"24",x"74",x"C3",x"05",x"90",x"D5",x"D2",x"31",x"4C",x"13",x"C4",x"94",x"6F",x"54",x"DA",x"94",x"A0",x"67",x"45",x"56",x"79",x"57",x"86",x"9A",x"3D",x"39",x"94",x"DD",x"BB",x"A8",x"BB",x"6D",x"D3",x"F4",x"A4",x"28",x"3A",x"75",x"4D",x"37",x"7C",x"02",x"5B",x"34",x"55",x"C3",x"B4",x"49",x"CC",x"59",x"E7",x"01",x"FF",
		x"60",x"AD",x"CF",x"85",x"3D",x"AA",x"E3",x"8E",x"A1",x"46",x"73",x"A9",x"5C",x"32",x"BA",x"5A",x"5C",x"D5",x"A3",x"75",x"E9",x"9A",x"4F",x"48",x"8F",x"C4",x"A0",x"80",x"B2",x"43",x"0D",x"D0",x"F5",x"A8",x"02",x"9A",x"2A",x"01",x"05",x"B4",x"EC",x"C6",x"80",x"52",x"8C",x"53",x"9E",x"32",x"7A",x"98",x"6D",x"1A",x"59",x"6E",x"14",x"A6",x"F1",x"78",x"A4",x"A9",x"88",x"87",x"E6",x"EC",x"91",x"E6",x"18",x"5E",x"EA",x"8B",x"46",x"12",x"AB",x"A6",x"C7",x"58",x"6D",x"51",x"8A",x"E1",x"11",x"69",x"3A",x"C4",x"39",x"BB",x"5B",x"4C",x"10",x"00",x"D1",x"79",x"E9",x"1A",x"9E",x"B5",x"C5",x"A0",x"55",x"64",x"AA",x"47",x"0A",x"43",x"30",x"1C",x"A6",x"15",x"7A",x"F4",x"39",x"6B",x"70",x"54",x"E5",x"35",x"D4",x"E4",x"C9",x"91",x"73",x"D6",x"50",x"73",x"24",x"47",x"CC",x"59",x"7D",x"2D",x"11",x"92",x"39",x"67",x"F5",x"2D",x"85",x"B1",x"D7",x"EC",x"D2",x"D4",x"20",x"8E",x"D1",x"55",x"19",x"90",x"90",x"84",x"02",x"56",x"14",x"1A",x"79",x"F3",x"EA",x"AC",x"59",x"7B",x"24",x"25",x"18",x"79",x"54",x"E7",x"92",x"B4",x"66",x"62",x"EA",x"A9",x"81",x"01",x"B1",x"7A",x"20",x"A0",x"CB",x"30",x"10",x"40",x"0A",x"14",x"2D",x"2D",x"A9",x"2C",x"C3",x"07",x"B7",x"28",x"55",x"2F",x"D7",x"0C",x"D3",x"82",x"DC",x"BC",x"CD",x"33",x"6A",x"73",x"53",x"F3",x"32",x"AF",x"A8",x"CD",x"49",x"C3",x"53",x"BD",x"A2",x"36",x"27",x"0E",x"4F",x"F5",x"9C",x"D2",x"DC",x"30",x"3C",x"CC",x"BD",x"66",x"F3",x"FC",x"90",x"72",x"F1",x"D9",x"25",x"F2",x"83",x"2B",x"C5",x"9A",x"94",x"32",x"4C",x"2A",x"F3",x"48",x"DE",x"DA",x"38",x"28",x"C2",x"23",x"59",x"1B",x"D3",x"A2",x"48",x"37",x"67",x"AD",x"4F",x"93",x"22",x"DC",x"93",x"3A",x"37",x"76",x"89",x"4C",x"8B",x"A2",x"BC",x"D0",x"A4",x"52",x"75",x"B6",x"08",x"43",x"A7",x"6C",x"D5",x"B6",x"AA",x"88",x"9D",x"32",x"55",x"5B",x"AB",x"36",x"0E",x"F6",x"16",x"5B",x"23",x"C6",x"34",x"31",x"8B",x"A3",x"35",x"1B",x"52",x"63",x"ED",x"B0",x"2C",x"0F",x"FF",
		x"60",x"23",x"EB",x"2E",x"83",x"C2",x"97",x"8C",x"B0",x"C6",x"10",x"F3",x"5A",x"32",x"FC",x"DA",x"C4",x"CD",x"A6",x"76",x"73",x"EB",x"AE",x"34",x"77",x"CB",x"06",x"A8",x"B1",x"D5",x"01",x"4B",x"4E",x"82",x"01",x"8A",x"31",x"1F",x"61",x"4D",x"A1",x"5A",x"D9",x"A6",x"F9",x"B5",x"AA",x"99",x"66",x"92",x"12",x"E4",x"8C",x"61",x"A1",x"AB",x"5A",x"90",x"0B",x"A6",x"45",x"CD",x"1A",x"61",x"CE",x"EC",x"96",x"B9",x"B8",x"A5",x"35",x"8B",x"A8",x"E7",x"6C",x"05",x"CC",x"51",x"61",x"80",x"D9",x"2A",x"0D",x"B0",x"46",x"07",x"03",x"D6",x"DD",x"60",x"C0",x"DA",x"E3",x"02",x"98",x"39",x"AD",x"85",x"C5",x"A9",x"69",x"65",x"ED",x"16",x"E6",x"18",x"11",x"9E",x"73",x"5A",x"18",x"4B",x"A7",x"85",x"CF",x"69",x"61",x"9A",x"19",x"1E",x"55",x"A5",x"45",x"B9",x"66",x"9A",x"75",x"5D",x"07",x"54",x"A7",x"45",x"80",x"E1",x"C5",x"08",x"10",x"94",x"A4",x"8B",x"72",x"32",x"8F",x"A8",x"2A",x"2E",x"4C",x"A5",x"D2",x"23",x"66",x"9B",x"30",x"CD",x"4C",x"8B",x"AA",x"AA",x"C2",x"DC",x"32",x"DC",x"BB",x"AA",x"00",x"72",x"15",x"1D",x"55",x"29",x"59",x"2A",x"5D",x"B6",x"95",x"A9",x"65",x"6A",x"D4",x"D4",x"51",x"65",x"37",x"69",x"EE",x"4B",x"46",x"93",x"62",x"A7",x"85",x"CF",x"69",x"6D",x"EC",x"AD",x"D6",x"D1",x"B8",x"F5",x"61",x"46",x"B8",x"D4",x"94",x"36",x"F8",x"E6",x"99",x"E4",x"73",x"DA",x"10",x"BA",x"A6",x"59",x"B8",x"2D",x"43",x"58",x"62",x"19",x"D6",x"74",x"4C",x"B1",x"A4",x"79",x"79",x"BD",x"31",x"A7",x"A2",x"96",x"A5",x"F1",x"CB",x"12",x"27",x"45",x"9B",x"AE",x"29",x"6B",x"9A",x"D8",x"A1",x"D5",x"24",x"2C",x"E9",x"62",x"A4",x"DB",x"2C",x"37",x"E6",x"45",x"99",x"6A",x"8D",x"DC",x"90",x"3A",x"5B",x"95",x"A6",x"56",x"53",x"6E",x"54",x"A9",x"D6",x"F8",x"01",x"FF",
		x"60",x"23",x"EA",x"AE",x"55",x"D3",x"D6",x"8C",x"B0",x"0D",x"E7",x"D4",x"98",x"23",x"80",x"52",x"CC",x"04",x"50",x"A7",x"99",x"02",x"BA",x"1F",x"15",x"C0",x"D2",x"A5",x"A0",x"80",x"EE",x"DA",x"04",x"D0",x"4A",x"4A",x"09",x"72",x"C7",x"70",x"F7",x"D6",x"2D",x"48",x"15",x"33",x"D4",x"17",x"8D",x"20",x"26",x"F1",x"0A",x"9F",x"35",x"C2",x"DC",x"CC",x"5C",x"63",x"F6",x"08",x"4B",x"E1",x"90",x"E8",x"B2",x"2D",x"6E",x"59",x"9C",x"3C",x"62",x"29",x"60",x"8E",x"29",x"03",x"CC",x"D5",x"E9",x"80",x"39",x"D3",x"1C",x"30",x"BA",x"89",x"02",x"46",x"75",x"6F",x"E1",x"18",x"61",x"66",x"96",x"76",x"A4",x"D9",x"AA",x"79",x"7B",x"E5",x"11",x"A7",x"EC",x"E1",x"51",x"53",x"46",x"9C",x"43",x"55",x"BA",x"2D",x"19",x"51",x"8E",x"15",x"69",x"31",x"67",x"A4",x"39",x"45",x"84",x"75",x"1D",x"97",x"D6",x"18",x"61",x"5C",x"69",x"14",x"30",x"44",x"27",x"03",x"52",x"10",x"37",x"71",x"4E",x"6E",x"E1",x"DD",x"C8",x"C5",x"C5",x"6E",x"A4",x"79",x"9B",x"10",x"15",x"33",x"91",x"EE",x"4D",x"18",x"30",x"44",x"27",x"03",x"16",x"8D",x"60",x"C0",x"F5",x"11",x"00",x"25",x"ED",x"D1",x"58",x"C5",x"62",x"8F",x"A4",x"57",x"13",x"34",x"9F",x"3B",x"E2",x"15",x"4C",x"41",x"7D",x"CD",x"88",x"46",x"0A",x"03",x"CD",x"D5",x"23",x"19",x"C1",x"18",x"AC",x"5B",x"8F",x"7C",x"5A",x"65",x"94",x"ED",x"34",x"CA",x"E1",x"8D",x"41",x"A6",x"D3",x"A8",x"67",x"70",x"01",x"A9",x"CE",x"A3",x"9B",x"29",x"15",x"24",x"3A",x"8F",x"7E",x"A6",x"34",x"D0",x"D8",x"3C",x"C6",x"51",x"5A",x"41",x"22",x"F3",x"98",x"66",x"6E",x"07",x"F2",x"CE",x"6D",x"EE",x"D1",x"18",x"AA",x"17",x"87",x"72",x"44",x"55",x"E2",x"5C",x"ED",x"9A",x"E1",x"8C",x"40",x"27",x"13",x"6A",x"67",x"0C",x"01",x"A9",x"4E",x"6E",x"6D",x"8A",x"85",x"A7",x"5A",x"87",x"B1",x"6A",x"51",x"DD",x"4C",x"24",x"A6",x"C4",x"D9",x"E2",x"CC",x"14",x"59",x"A3",x"62",x"AF",x"25",x"CB",x"0F",x"FF",
		x"60",x"23",x"19",x"D9",x"8B",x"DD",x"96",x"AE",x"B8",x"27",x"0F",x"71",x"9F",x"3B",x"A2",x"56",x"53",x"24",x"75",x"A9",x"0B",x"5A",x"15",x"B6",x"8C",x"9A",x"0E",x"A8",x"DD",x"2D",x"00",x"CD",x"A7",x"28",x"60",x"9B",x"51",x"50",x"40",x"0D",x"12",x"23",x"EA",x"B5",x"4C",x"CD",x"D2",x"B4",x"20",x"77",x"72",x"35",x"6D",x"D2",x"FC",x"98",x"45",x"23",x"E5",x"D1",x"08",x"52",x"08",x"CB",x"90",x"45",x"23",x"4C",x"BE",x"D4",x"CA",x"16",x"8D",x"38",x"05",x"8F",x"B0",x"1C",x"AD",x"80",x"64",x"5D",x"05",x"90",x"AD",x"99",x"00",x"82",x"55",x"35",x"41",x"0E",x"21",x"66",x"9E",x"D4",x"F9",x"D9",x"B9",x"45",x"5A",x"BD",x"10",x"66",x"57",x"E6",x"61",x"AB",x"09",x"90",x"5D",x"F8",x"70",x"93",x"9F",x"74",x"93",x"45",x"C3",x"CD",x"B1",x"C2",x"3D",x"E6",x"0C",x"A7",x"44",x"F3",x"C8",x"9A",x"3A",x"EC",x"96",x"58",x"23",x"27",x"EA",x"70",x"9A",x"62",x"9A",x"EE",x"38",x"C5",x"1E",x"91",x"28",x"73",x"63",x"01",x"01",x"92",x"9F",x"70",x"4E",x"8E",x"95",x"EE",x"3E",x"C7",x"B8",x"25",x"79",x"78",x"D4",x"54",x"67",x"B7",x"28",x"92",x"D1",x"55",x"99",x"D3",x"14",x"49",x"77",x"DB",x"11",x"40",x"D1",x"E6",x"0A",x"70",x"42",x"62",x"E4",x"39",x"4E",x"A6",x"64",x"95",x"56",x"C6",x"96",x"A9",x"D9",x"55",x"46",x"51",x"5C",x"B5",x"B9",x"2D",x"19",x"55",x"31",x"D5",x"1E",x"BA",x"64",x"34",x"D9",x"4C",x"7B",x"F0",x"9A",x"D6",x"86",x"3C",x"15",x"AE",x"AB",x"5B",x"1B",x"52",x"54",x"1B",x"37",x"69",x"5D",x"28",x"E1",x"65",x"D4",x"A4",x"0D",x"B1",x"A4",x"56",x"61",x"DB",x"36",x"A4",x"1A",x"9A",x"69",x"F6",x"DB",x"98",x"5A",x"98",x"97",x"DA",x"6B",x"53",x"AE",x"29",x"3A",x"12",x"AF",x"CD",x"B9",x"85",x"D8",x"52",x"D2",x"B2",x"A4",x"6E",x"E2",x"43",x"4D",x"42",x"97",x"16",x"6B",x"16",x"AF",x"0E",x"43",x"BE",x"14",x"A9",x"B2",x"C5",x"AD",x"F9",x"8A",x"B7",x"F2",x"1C",x"B7",x"E7",x"25",x"D6",x"4E",x"4D",x"DC",x"54",x"26",x"5B",x"06",x"37",x"51",x"73",x"6C",x"58",x"ED",x"3A",x"5A",x"2C",x"A1",x"51",x"95",x"6B",x"65",x"B2",x"85",x"86",x"D9",x"61",x"B1",x"1F",x"FF",
		x"60",x"C6",x"4D",x"19",x"D3",x"A3",x"4C",x"25",x"33",x"24",x"89",x"1C",x"B3",x"54",x"B4",x"98",x"29",x"62",x"BC",x"50",x"53",x"53",x"A2",x"B4",x"CE",x"22",x"4D",x"CB",x"89",x"52",x"32",x"86",x"34",x"2D",x"27",x"76",x"29",x"3B",x"5C",x"8C",x"9C",x"29",x"A5",x"62",x"74",x"71",x"72",x"A1",x"E6",x"AE",x"D1",x"C5",x"CD",x"95",x"4A",x"2A",x"27",x"17",x"2F",x"37",x"4A",x"C9",x"98",x"5C",x"C2",x"9C",x"28",x"3D",x"B5",x"62",x"CA",x"EB",x"D2",x"10",x"C7",x"C9",x"AE",x"A9",x"53",x"82",x"83",x"6A",x"B1",x"BE",x"6E",x"09",x"09",x"89",x"F5",x"00",x"FF",
		x"60",x"4E",x"09",x"91",x"32",x"3B",x"42",x"26",x"D5",x"47",x"9D",x"4C",x"AB",x"D2",x"64",x"57",x"B4",x"B2",x"3C",x"76",x"93",x"7C",x"92",x"AA",x"CE",x"8A",x"4D",x"F4",x"51",x"3B",x"CB",x"22",x"17",x"D1",x"67",x"AD",x"18",x"8F",x"5C",x"A4",x"50",x"38",x"73",x"AC",x"4A",x"D1",x"62",x"E6",x"8C",x"D6",x"22",x"C5",x"49",x"99",x"DA",x"AA",x"4A",x"97",x"20",x"57",x"0A",x"4B",x"1F",x"5D",x"E2",x"3C",x"29",x"34",x"BC",x"4C",x"29",x"72",x"63",x"B3",x"D6",x"5A",x"A9",x"CD",x"49",x"D4",x"96",x"4B",x"85",x"BE",x"54",x"56",x"49",x"69",x"E4",x"86",x"52",x"C8",x"35",x"B5",x"A6",x"18",x"CB",x"10",x"15",x"F7",x"C4",x"0F",x"FF",
		x"60",x"4A",x"2F",x"C9",x"55",x"D5",x"12",x"17",x"2D",x"27",x"0A",x"2B",x"6F",x"D0",x"D4",x"94",x"A9",x"24",x"33",x"76",x"53",x"73",x"C2",x"A1",x"A9",x"D8",x"4D",x"4B",x"19",x"4B",x"3B",x"2A",x"37",x"2D",x"06",x"2E",x"1F",x"6D",x"50",x"AC",x"9C",x"B0",x"B5",x"A2",x"42",x"73",x"4B",x"C3",x"A2",x"8A",x"4A",x"25",x"AC",x"83",x"82",x"42",x"67",x"86",x"B4",x"0E",x"72",x"71",x"AE",x"19",x"CA",x"3A",x"D9",x"D9",x"35",x"A6",x"2B",x"EB",x"64",x"27",x"95",x"56",x"21",x"AB",x"0D",x"83",x"CB",x"6A",x"BA",x"AA",x"24",x"28",x"ED",x"AC",x"69",x"FA",x"3A",x"D0",x"C4",x"22",x"26",x"02",x"DA",x"B1",x"44",x"40",x"9B",x"9E",x"08",x"68",x"DB",x"E2",x"01",x"FF",
		x"60",x"25",x"69",x"DA",x"D4",x"C4",x"56",x"8F",x"28",x"45",x"49",x"F6",x"5E",x"32",x"A2",x"14",x"23",x"95",x"72",x"CD",x"08",x"A2",x"CE",x"2E",x"B2",x"34",x"C3",x"0B",x"B6",x"DA",x"20",x"9C",x"34",x"C7",x"BA",x"68",x"93",x"70",x"E3",x"1C",x"6B",x"AC",x"85",x"32",x"0E",x"08",x"A0",x"69",x"0B",x"05",x"34",x"99",x"69",x"80",x"69",x"55",x"0C",x"B0",x"52",x"AA",x"02",x"56",x"2C",x"13",x"C0",x"28",x"93",x"C5",x"AE",x"39",x"9D",x"58",x"E3",x"34",x"37",x"7B",x"36",x"77",x"6E",x"9B",x"DC",x"E4",x"C8",x"3D",x"24",x"9D",x"F3",x"AA",x"34",x"57",x"E1",x"B4",x"0C",x"E8",x"9C",x"49",x"01",x"3D",x"98",x"26",x"BF",x"B7",x"0E",x"21",x"72",x"D2",x"E2",x"12",x"85",x"3C",x"A5",x"6B",x"8B",x"83",x"37",x"CB",x"E4",x"D5",x"2D",x"F5",x"29",x"35",x"83",x"16",x"B7",x"CC",x"D7",x"D4",x"4C",x"5C",x"5C",x"72",x"3F",x"38",x"53",x"65",x"71",x"6A",x"53",x"8C",x"30",x"37",x"BB",x"02",x"28",x"C1",x"55",x"00",x"C3",x"75",x"B8",x"B8",x"9B",x"30",x"35",x"77",x"A2",x"92",x"AC",x"C2",x"C3",x"DD",x"8E",x"C9",x"8A",x"F4",x"A8",x"70",x"AB",x"0C",x"68",x"26",x"3C",x"85",x"61",x"73",x"84",x"AB",x"D3",x"12",x"84",x"4E",x"ED",x"29",x"9D",x"5A",x"10",x"33",x"97",x"45",x"34",x"1E",x"61",x"8E",x"66",x"66",x"B1",x"78",x"44",x"39",x"AA",x"79",x"56",x"ED",x"91",x"E4",x"24",x"61",x"D5",x"51",x"46",x"56",x"63",x"A8",x"49",x"D5",x"19",x"45",x"89",x"21",x"66",x"53",x"A5",x"55",x"C9",x"84",x"26",x"67",x"D4",x"D6",x"26",x"A7",x"1E",x"5A",x"6A",x"5A",x"57",x"82",x"99",x"72",x"26",x"6A",x"7D",x"31",x"1A",x"26",x"ED",x"A8",x"74",x"C5",x"69",x"B0",x"B5",x"ED",x"32",x"D6",x"E8",x"A6",x"5C",x"B1",x"CB",x"5C",x"7D",x"88",x"C9",x"44",x"76",x"6B",x"92",x"62",x"C9",x"15",x"D9",x"AC",x"91",x"AB",x"95",x"54",x"64",x"02",x"30",x"1D",x"21",x"80",x"04",x"DC",x"05",x"90",x"A1",x"BA",x"00",x"3A",x"54",x"23",x"80",x"35",x"66",x"08",x"90",x"D1",x"3D",x"4D",x"31",x"55",x"93",x"F6",x"9C",x"36",x"25",x"DF",x"AD",x"6C",x"53",x"C7",x"94",x"75",x"B7",x"A9",x"CE",x"1D",x"53",x"72",x"9B",x"AC",x"31",x"B5",x"2C",x"59",x"97",x"1B",x"DB",x"9C",x"30",x"17",x"29",x"6E",x"E8",x"6D",x"CC",x"1C",x"B9",x"9B",x"4B",x"B4",x"32",x"6B",x"74",x"99",x"C2",x"6E",x"D9",x"AD",x"31",x"BA",x"B3",x"59",x"E4",x"36",x"35",x"67",x"21",x"AA",x"B3",x"C6",x"DC",x"AD",x"B9",x"A8",x"6D",x"1A",x"4B",x"B3",x"EE",x"86",x"BE",x"39",x"AD",x"D5",x"9A",x"2B",x"F4",x"1A",x"06",x"0C",x"E8",x"C2",x"80",x"49",x"5D",x"05",x"70",x"45",x"98",x"00",x"36",x"11",x"0B",x"63",x"35",x"E6",x"CA",x"D1",x"D0",x"4D",x"91",x"96",x"A5",x"46",x"69",x"37",x"07",x"76",x"C6",x"6E",x"4B",x"D2",x"1C",x"F5",x"38",x"7B",x"CD",x"2D",x"53",x"8A",x"15",x"6C",x"3B",x"B5",x"4D",x"D9",x"75",x"AA",x"D4",x"D5",x"32",x"A7",x"5C",x"A6",x"3E",x"E3",x"CA",x"92",x"42",x"BB",x"92",x"5F",x"31",x"4B",x"0A",x"25",x"2C",x"5E",x"3B",x"AC",x"3E",x"4E",x"88",x"D4",x"D5",x"B0",x"FA",x"BC",x"CA",x"5E",x"63",x"DC",x"E6",x"DB",x"88",x"58",x"4F",x"35",x"BB",x"2B",x"C7",x"1C",x"39",x"45",x"6D",x"B6",x"6E",x"88",x"64",x"9C",x"07",x"FF",
		x"60",x"A9",x"6A",x"5E",x"98",x"32",x"1B",x"B7",x"AC",x"64",x"16",x"37",x"DD",x"D2",x"92",x"98",x"38",x"43",x"75",x"75",x"4B",x"62",x"75",x"29",x"A3",x"D5",x"25",x"8D",x"93",x"AD",x"59",x"16",x"97",x"24",x"2D",x"B2",x"66",x"59",x"9C",x"B2",x"F2",x"A8",x"84",x"6C",x"8E",x"02",x"C6",x"98",x"56",x"C0",x"6C",x"A5",x"0A",x"58",x"7D",x"5D",x"01",x"A3",x"97",x"2B",x"A0",x"6F",x"8B",x"11",x"A5",x"CA",x"69",x"D1",x"51",x"47",x"9C",x"72",x"86",x"BB",x"CF",x"19",x"49",x"4A",x"1D",x"EE",x"B6",x"64",x"44",x"A9",x"74",x"98",x"C7",x"E2",x"11",x"C6",x"96",x"E6",x"55",x"75",x"5A",x"90",x"93",x"87",x"FA",x"54",x"05",x"01",x"A4",x"C2",x"8E",x"80",x"6C",x"36",x"15",x"50",x"E5",x"A6",x"02",x"AA",x"9A",x"60",x"40",x"A3",x"EE",x"08",x"E8",x"32",x"8C",x"15",x"9E",x"95",x"BB",x"B9",x"ED",x"92",x"B5",x"1C",x"C1",x"9C",x"51",x"47",x"5A",x"9B",x"07",x"47",x"C6",x"1D",x"69",x"AD",x"5E",x"EA",x"55",x"67",x"24",x"A5",x"45",x"99",x"65",x"9D",x"16",x"E7",x"12",x"69",x"5E",x"75",x"5B",x"98",x"52",x"A5",x"59",x"4E",x"69",x"61",x"0C",x"5D",x"A6",x"31",x"BB",x"05",x"21",x"75",x"AA",x"79",x"DD",x"E6",x"87",x"90",x"E5",x"6E",x"E1",x"5A",x"10",x"83",x"66",x"44",x"86",x"6D",x"49",x"29",x"1E",x"A6",x"11",x"BA",x"E4",x"25",x"55",x"78",x"78",x"D9",x"94",x"E7",x"5C",x"69",x"1E",x"55",x"4B",x"98",x"52",x"86",x"65",x"54",x"4D",x"59",x"4C",x"E9",x"16",x"1E",x"35",x"25",x"B1",x"B2",x"65",x"59",x"B4",x"94",x"E4",x"83",x"56",x"C6",x"4B",x"53",x"9C",x"27",x"64",x"69",x"2C",x"4A",x"51",x"9E",x"90",x"A5",x"31",x"2B",x"85",x"E5",x"42",x"BA",x"44",x"2D",x"13",x"D6",x"4B",x"6E",x"62",x"1D",x"01",x"01",x"D5",x"57",x"84",x"A8",x"74",x"D6",x"08",x"4F",x"37",x"DA",x"5C",x"24",x"BC",x"AB",x"CA",x"A8",x"72",x"F1",x"B0",x"EC",x"38",x"A3",x"C8",x"21",x"42",x"7D",x"E2",x"BA",x"2A",x"7B",x"75",x"95",x"B2",x"EB",x"52",x"A7",x"C3",x"CD",x"BC",x"CA",x"48",x"8B",x"49",x"35",x"F6",x"29",x"23",x"CD",x"49",x"D4",x"4D",x"57",x"97",x"34",x"55",x"B2",x"0C",x"D9",x"9C",x"B2",x"58",x"D9",x"2D",x"5D",x"99",x"2B",x"72",x"88",x"30",x"9F",x"2A",x"C0",x"00",x"A8",x"3C",x"43",x"9A",x"6D",x"A8",x"58",x"24",x"4B",x"89",x"0F",x"A5",x"15",x"21",x"AD",x"C5",x"51",x"5D",x"AA",x"F8",x"94",x"91",x"24",x"39",x"69",x"16",x"93",x"47",x"96",x"A3",x"87",x"59",x"37",x"19",x"45",x"CD",x"AE",x"EA",x"39",x"67",x"54",x"AD",x"84",x"88",x"C7",x"DC",x"D1",x"B4",x"9E",x"2C",x"E6",x"6B",x"46",x"D7",x"52",x"91",x"A4",x"AD",x"69",x"43",x"CD",x"8E",x"DE",x"BA",x"B9",x"8D",x"A5",x"36",x"6B",x"61",x"97",x"36",x"95",x"5E",x"A4",x"85",x"5D",x"DB",x"9C",x"4B",x"90",x"B6",x"B4",x"2B",x"4B",x"A9",x"C6",x"5A",x"DA",x"2E",x"6C",x"35",x"3A",x"4B",x"78",x"DD",x"70",x"D4",x"50",x"CC",x"E5",x"DD",x"08",x"90",x"4D",x"92",x"04",x"18",x"90",x"5C",x"22",x"01",x"62",x"70",x"42",x"40",x"F0",x"4E",x"0F",x"FF",
		x"60",x"0C",x"98",x"96",x"51",x"00",x"33",x"08",x"09",x"60",x"34",x"D1",x"16",x"F5",x"E6",x"A6",x"22",x"C9",x"5A",x"12",x"B3",x"69",x"64",x"57",x"6E",x"69",x"B6",x"13",x"C9",x"FE",x"B8",x"65",x"D9",x"4C",x"A4",x"FA",x"ED",x"96",x"66",x"BF",x"1E",x"96",x"53",x"42",x"12",x"53",x"A4",x"C5",x"44",x"61",x"40",x"96",x"5C",x"04",x"68",x"1E",x"CD",x"C5",x"31",x"BA",x"46",x"55",x"E5",x"92",x"66",x"DB",x"91",x"12",x"73",x"5A",x"96",x"CD",x"44",x"AA",x"D5",x"6E",x"51",x"8C",x"66",x"6A",x"3B",x"A6",x"25",x"DE",x"46",x"BA",x"47",x"23",x"53",x"64",x"63",x"A6",x"6A",x"76",x"11",x"10",x"A5",x"29",x"02",x"A2",x"36",x"43",x"40",x"D6",x"AE",x"08",x"B0",x"5C",x"3D",x"84",x"C9",x"86",x"5A",x"54",x"93",x"14",x"47",x"6F",x"6E",x"6E",x"B1",x"4B",x"1C",x"82",x"96",x"88",x"AF",x"6A",x"99",x"8F",x"EE",x"8E",x"DD",x"B9",x"E5",x"CE",x"A5",x"27",x"55",x"E7",x"56",x"06",x"1B",x"96",x"E8",x"7D",x"5B",x"13",x"79",x"59",x"91",x"F9",x"6B",x"6D",x"D4",x"E1",x"41",x"E2",x"AF",x"75",x"51",x"A4",x"15",x"AB",x"BF",x"D6",x"67",x"E5",x"5E",x"22",x"FA",x"DA",x"98",x"54",x"78",x"31",x"FB",x"2F",x"53",x"14",x"EE",x"A9",x"AA",x"AF",x"4C",x"C1",x"78",x"04",x"6B",x"BE",x"34",x"47",x"65",x"E1",x"C6",x"FA",x"CB",x"12",x"B5",x"85",x"19",x"E7",x"2B",x"4B",x"36",x"62",x"1A",x"EA",x"2F",x"CC",x"39",x"08",x"99",x"87",x"6D",x"B2",x"24",x"E9",x"56",x"2C",x"5A",x"DD",x"DA",x"AD",x"96",x"84",x"4B",x"56",x"73",x"55",x"1C",x"6E",x"1E",x"85",x"AD",x"59",x"A8",x"BB",x"BB",x"92",x"07",x"FF",
		x"60",x"08",x"A8",x"2E",x"83",x"00",x"2D",x"44",x"10",x"A0",x"C5",x"F4",x"50",x"05",x"9F",x"A5",x"1A",x"4E",x"53",x"E5",x"77",x"98",x"D4",x"5A",x"69",x"55",x"8C",x"35",x"50",x"9D",x"78",x"54",x"C5",x"C4",x"8A",x"74",x"93",x"51",x"35",x"AD",x"93",x"1C",x"4D",x"46",x"59",x"75",x"B4",x"4B",x"D6",x"19",x"45",x"31",x"19",x"9A",x"59",x"67",x"14",x"C5",x"58",x"58",x"65",x"E5",x"91",x"B7",x"E0",x"C6",x"E1",x"B3",x"47",x"DE",x"B2",x"AA",x"44",x"4E",x"19",x"79",x"0F",x"CA",x"E2",x"55",x"65",x"64",x"C3",x"09",x"5B",x"44",x"D8",x"91",x"34",x"63",x"E2",x"EE",x"61",x"5B",x"9C",x"AD",x"B9",x"A9",x"C7",x"6A",x"71",x"31",x"6A",x"EE",x"51",x"AB",x"E5",x"D5",x"89",x"69",x"F8",x"A4",x"52",x"D4",x"C0",x"CA",x"19",x"65",x"42",x"DE",x"BD",x"B0",x"44",x"56",x"19",x"45",x"F5",x"A1",x"4A",x"51",x"77",x"D4",x"45",x"97",x"B8",x"F6",x"9D",x"D1",x"D6",x"A0",x"A1",x"32",x"4D",x"C6",x"D0",x"B5",x"68",x"59",x"D5",x"6E",x"73",x"0F",x"AE",x"EA",x"1D",x"32",x"2D",x"CB",x"BA",x"A8",x"79",x"14",x"02",x"74",x"81",x"C1",x"80",x"21",x"45",x"47",x"5E",x"B5",x"A9",x"59",x"A4",x"1D",x"49",x"8F",x"2A",x"E4",x"D5",x"64",x"C4",x"C5",x"88",x"78",x"4E",x"95",x"96",x"64",x"23",x"EA",x"D9",x"91",x"55",x"96",x"85",x"AA",x"78",x"47",x"72",x"51",x"E4",x"96",x"61",x"29",x"3B",x"05",x"5E",x"69",x"AB",x"A5",x"E5",x"10",x"58",x"6D",x"E5",x"1E",x"76",x"52",x"18",x"15",x"65",x"74",x"88",x"49",x"51",x"52",x"62",x"95",x"65",x"D8",x"25",x"25",x"A8",x"68",x"74",x"14",x"00",x"02",x"10",x"5D",x"52",x"A2",x"10",x"26",x"D8",x"6D",x"72",x"8B",x"83",x"ED",x"32",x"D1",x"45",x"25",x"76",x"A1",x"8B",x"D5",x"16",x"B5",x"D8",x"BB",x"6C",x"61",x"DB",x"D2",x"D2",x"68",x"BD",x"59",x"AC",x"73",x"CA",x"83",x"33",x"57",x"8D",x"D6",x"02",x"68",x"BD",x"5A",x"00",x"7D",x"4C",x"09",x"A0",x"8F",x"8A",x"52",x"D5",x"C8",x"A6",x"19",x"4D",x"5A",x"53",x"0D",x"9B",x"45",x"34",x"6D",x"43",x"53",x"61",x"14",x"31",x"3B",x"4C",x"25",x"B0",x"88",x"79",x"DC",x"30",x"D7",x"A2",x"C2",x"6A",x"49",x"DD",x"9A",x"23",x"9B",x"79",x"D8",x"36",x"7B",x"76",x"EC",x"96",x"19",x"9B",x"1D",x"D9",x"B0",x"6B",x"55",x"E3",x"07",x"FF",
		x"60",x"0C",x"A8",x"5C",x"93",x"01",x"95",x"9B",x"85",x"32",x"33",x"AB",x"52",x"8B",x"DD",x"F2",x"10",x"3B",x"54",x"BB",x"CA",x"28",x"B2",x"89",x"34",x"A9",x"B9",x"23",x"6F",x"DE",x"45",x"AD",x"96",x"8C",x"AC",x"87",x"14",x"96",x"5C",x"3D",x"B2",x"E6",x"54",x"B8",x"6A",x"75",x"4B",x"6B",x"54",x"B2",x"CE",x"CE",x"2D",x"29",x"49",x"28",x"3B",x"DA",x"B4",x"B8",x"34",x"96",x"92",x"58",x"DD",x"A2",x"DC",x"84",x"DB",x"B4",x"4B",x"8B",x"73",x"13",x"4E",x"B7",x"B4",x"2D",x"C9",x"55",x"D9",x"C3",x"D3",x"B6",x"34",x"45",x"13",x"8D",x"E8",x"5A",x"D2",x"A2",x"CD",x"24",x"BC",x"99",x"00",x"BA",x"4D",x"11",x"40",x"37",x"C3",x"02",x"68",x"66",x"14",x"18",x"90",x"87",x"B0",x"00",x"5A",x"2E",x"6B",x"59",x"F5",x"6A",x"A6",x"59",x"7B",x"14",x"25",x"49",x"48",x"55",x"9C",x"50",x"44",x"25",x"5E",x"9A",x"91",x"43",x"9E",x"35",x"5B",x"4A",x"45",x"76",x"79",x"32",x"1C",x"6A",x"1D",x"A5",x"65",x"35",x"7B",x"B0",x"65",x"95",x"91",x"D5",x"E2",x"C5",x"19",x"55",x"46",x"5A",x"8A",x"A7",x"44",x"56",x"19",x"49",x"CE",x"19",x"6A",x"55",x"75",x"C4",x"29",x"B7",x"AB",x"67",x"D5",x"11",x"A5",x"D8",x"A1",x"96",x"53",x"46",x"14",x"42",x"A7",x"69",x"4E",x"19",x"91",x"CF",x"99",x"6A",x"15",x"B7",x"45",x"3E",x"66",x"9A",x"85",x"B5",x"92",x"C4",x"18",x"61",x"96",x"62",x"48",x"9C",x"4B",x"84",x"58",x"86",x"49",x"71",x"4A",x"ED",x"6A",x"51",x"A6",x"E4",x"29",x"B4",x"A9",x"59",x"95",x"91",x"06",x"53",x"EE",x"2E",x"8B",x"47",x"16",x"6D",x"96",x"B3",x"2C",x"19",x"59",x"F0",x"D5",x"4A",x"BA",x"78",x"A4",x"C1",x"55",x"2B",x"E9",x"E2",x"96",x"F9",x"D0",x"25",x"68",x"8B",x"53",x"6A",x"73",x"37",x"53",x"4C",x"09",x"A9",x"AB",x"53",x"C2",x"31",x"B5",x"0C",x"7E",x"4C",x"0A",x"47",x"D3",x"D2",x"F9",x"DE",x"25",x"5C",x"73",x"4A",x"19",x"5A",x"17",x"4B",x"57",x"69",x"79",x"E8",x"59",x"94",x"1D",x"B7",x"E5",x"A1",x"54",x"B3",x"77",x"9D",x"56",x"84",x"96",x"29",x"36",x"51",x"53",x"1A",x"F2",x"9A",x"7B",x"94",x"21",x"40",x"B6",x"A1",x"04",x"C8",x"3A",x"13",x"03",x"0C",x"C8",x"7C",x"93",x"01",x"83",x"85",x"70",x"80",x"00",x"83",x"87",x"51",x"00",x"18",x"90",x"8B",x"89",x"CB",x"73",x"0A",x"52",x"F7",x"24",x"A1",x"8C",x"45",x"A8",x"5D",x"D3",x"A6",x"32",x"35",x"E2",x"36",x"E9",x"52",x"AA",x"D2",x"D0",x"C2",x"A2",x"71",x"A9",x"6B",x"45",x"D3",x"8A",x"5A",x"AD",x"A9",x"91",x"D4",x"3A",x"23",x"B7",x"AE",x"19",x"61",x"ED",x"0C",x"D5",x"FA",x"21",x"55",x"B4",x"33",x"52",x"1B",x"A7",x"35",x"A6",x"CC",x"4A",x"6D",x"5A",x"C6",x"98",x"32",x"63",x"B7",x"65",x"59",x"57",x"72",x"4D",x"5A",x"B6",x"AE",x"43",x"D1",x"AC",x"4E",x"D8",x"B3",x"23",x"8E",x"8C",x"C8",x"E1",x"2C",x"9A",x"D9",x"2A",x"AC",x"B8",x"AB",x"0B",x"11",x"4B",x"8F",x"AC",x"EF",x"07",x"FF",
		x"60",x"A9",x"6A",x"99",x"85",x"34",x"EA",x"8C",x"62",x"96",x"0C",x"40",x"6D",x"3A",x"AA",x"D5",x"32",x"08",x"A9",x"ED",x"A8",x"67",x"29",x"07",x"92",x"76",x"AD",x"6E",x"41",x"58",x"52",x"B2",x"85",x"3A",x"48",x"8B",x"08",x"F4",x"E6",x"6A",x"6F",x"33",x"5C",x"C5",x"71",x"A8",x"83",x"F1",x"2C",x"61",x"DB",x"A5",x"4E",x"42",x"3B",x"D3",x"C8",x"8C",x"BA",x"08",x"9D",x"72",x"A6",x"37",x"AA",x"66",x"34",x"23",x"44",x"DB",x"A8",x"AA",x"B3",x"B0",x"D0",x"AE",x"A3",x"AA",x"49",x"CD",x"DC",x"BA",x"8C",x"B2",x"65",x"55",x"73",x"5F",x"3D",x"CA",x"96",x"55",x"D4",x"73",x"F5",x"28",x"5B",x"51",x"D5",x"C8",x"D6",x"A3",x"6A",x"45",x"55",x"3D",x"5B",x"8F",x"AA",x"16",x"55",x"F7",x"6A",x"33",x"EA",x"5A",x"54",x"52",x"7B",x"C9",x"68",x"4A",x"32",x"4E",x"8F",x"55",x"A3",x"29",x"49",x"39",x"C3",x"57",x"8D",x"B6",x"54",x"95",x"74",x"DB",x"DC",x"BA",x"52",x"C9",x"23",x"6D",x"75",x"EB",x"72",x"23",x"8F",x"F0",x"2C",x"AD",x"4F",x"55",x"34",x"34",x"D3",x"96",x"3E",x"17",x"76",x"97",x"68",x"9B",x"C6",x"92",x"4D",x"22",x"BC",x"75",x"E8",x"4B",x"31",x"CE",x"B0",x"CD",x"A9",x"2B",x"D9",x"C5",x"D2",x"BD",x"B6",x"B6",x"14",x"57",x"D1",x"8E",x"3B",x"CA",x"1A",x"24",x"C8",x"B7",x"F6",x"A8",x"9A",x"37",x"67",x"F5",x"39",x"AE",x"CB",x"89",x"CD",x"CC",x"DB",x"8A",x"2E",x"49",x"17",x"D7",x"A8",x"0D",x"04",x"A8",x"D2",x"A9",x"65",x"23",x"85",x"22",x"DB",x"DC",x"91",x"CC",x"10",x"02",x"9A",x"71",x"5B",x"B4",x"AC",x"09",x"49",x"BA",x"6D",x"E1",x"32",x"4A",x"EC",x"6B",x"79",x"44",x"CB",x"3B",x"8A",x"6F",x"A5",x"91",x"F4",x"68",x"64",x"16",x"4D",x"52",x"56",x"1D",x"5A",x"53",x"DA",x"0D",x"79",x"31",x"68",x"C5",x"99",x"64",x"54",x"C5",x"A9",x"3B",x"7B",x"E3",x"D1",x"94",x"E0",x"21",x"12",x"8D",x"47",x"57",x"43",x"84",x"51",x"34",x"19",x"7D",x"8D",x"E5",x"4A",x"D1",x"66",x"F4",x"CD",x"87",x"29",x"65",x"93",x"32",x"36",x"93",x"62",x"E8",x"8D",x"C3",x"58",x"2D",x"BB",x"70",x"39",x"49",x"53",x"75",x"EA",x"8A",x"E9",x"24",x"2D",x"25",x"78",x"30",x"55",x"92",x"32",x"57",x"EF",x"A1",x"98",x"49",x"D2",x"52",x"63",x"BA",x"60",x"26",x"09",x"6B",x"F5",x"66",x"42",x"59",x"C7",x"AD",x"D9",x"06",x"9B",x"7A",x"63",x"04",x"70",x"2F",x"49",x"00",x"4F",x"52",x"09",x"30",x"A0",x"19",x"01",x"06",x"36",x"45",x"C0",x"24",x"21",x"08",x"98",x"AC",x"EC",x"01",x"FF",
		x"60",x"0C",x"18",x"9A",x"55",x"01",x"2B",x"A5",x"08",x"60",x"EE",x"B4",x"94",x"65",x"4F",x"96",x"99",x"B5",x"5B",x"95",x"83",x"46",x"78",x"2C",x"69",x"5D",x"8E",x"51",x"AE",x"BE",x"A4",x"B5",x"39",x"56",x"73",x"C6",x"9C",x"56",x"E7",x"50",x"A3",x"1A",x"4B",x"52",x"95",x"43",x"A7",x"6B",x"DC",x"21",x"80",x"6F",x"66",x"08",x"F0",x"59",x"03",x"10",x"10",x"7A",x"04",x"01",x"62",x"8F",x"1C",x"4E",x"72",x"21",x"AE",x"5D",x"79",x"38",x"C9",x"69",x"B9",x"74",x"95",x"E4",x"86",x"E4",x"6E",x"92",x"55",x"01",x"80",x"01",x"C5",x"A5",x"11",x"40",x"A6",x"88",x"64",x"F8",x"D8",x"A1",x"A2",x"65",x"8A",x"16",x"7A",x"38",x"FB",x"04",x"2D",x"6A",x"08",x"1B",x"A2",x"36",x"A6",x"28",x"A1",x"B4",x"89",x"FA",x"D4",x"A2",x"F8",x"9C",x"2E",x"56",x"53",x"8B",x"E8",x"7D",x"A4",x"49",x"2C",x"4A",x"72",x"72",x"54",x"AA",x"51",x"53",x"01",x"AD",x"A8",x"2B",x"A0",x"25",x"33",x"A3",x"36",x"27",x"59",x"E1",x"52",x"8C",x"52",x"8D",x"5A",x"44",x"C4",x"2E",x"69",x"8D",x"64",x"E6",x"D1",x"A4",x"E5",x"29",x"B2",x"59",x"E6",x"E2",x"51",x"56",x"93",x"46",x"19",x"4D",x"47",x"3F",x"94",x"27",x"99",x"AE",x"0D",x"73",x"15",x"A2",x"EE",x"5A",x"C7",x"CD",x"55",x"91",x"86",x"7A",x"1D",x"B7",x"36",x"83",x"E6",x"E6",x"71",x"DD",x"96",x"AC",x"98",x"46",x"37",x"09",x"6B",x"31",x"A1",x"54",x"D9",x"E4",x"01",x"FF",
		x"60",x"21",x"1D",x"81",x"0D",x"D4",x"1B",x"A7",x"A0",x"05",x"15",x"90",x"4A",x"D5",x"DC",x"DA",x"84",x"49",x"22",x"F5",x"30",x"4B",x"21",x"31",x"F6",x"96",x"4D",x"CB",x"96",x"3C",x"95",x"1B",x"35",x"35",x"79",x"4B",x"21",x"6D",x"54",x"B4",x"E0",x"2C",x"59",x"32",x"56",x"D1",x"A3",x"55",x"33",x"C9",x"2A",x"C5",x"2E",x"26",x"94",x"D9",x"1B",x"1B",x"20",x"51",x"B3",x"62",x"0D",x"53",x"0E",x"62",x"6E",x"8D",x"91",x"1D",x"5B",x"A8",x"34",x"32",x"56",x"74",x"16",x"C6",x"D6",x"D8",x"05",x"C1",x"72",x"A9",x"46",x"EC",x"E1",x"65",x"EF",x"1A",x"E9",x"63",x"86",x"53",x"92",x"B8",x"67",x"97",x"1D",x"66",x"4E",x"1A",x"91",x"13",x"66",x"18",x"25",x"6B",x"58",x"4D",x"98",x"61",x"96",x"28",x"E1",x"DD",x"51",x"87",x"5D",x"9C",x"84",x"CE",x"D8",x"0E",x"5E",x"36",x"69",x"9A",x"5E",x"87",x"01",x"53",x"96",x"8F",x"B4",x"3A",x"0B",x"8D",x"8A",x"3C",x"F2",x"9A",x"55",x"25",x"B2",x"CC",x"68",x"5B",x"35",x"36",x"8F",x"46",x"BA",x"15",x"40",x"71",x"E2",x"00",x"00",x"0C",x"C8",x"96",x"CD",x"85",x"3D",x"B8",x"B2",x"68",x"A3",x"94",x"E4",x"20",x"A6",x"9A",x"73",x"58",x"1E",x"B5",x"A9",x"BA",x"37",x"02",x"20",x"40",x"53",x"6C",x"0C",x"18",x"9A",x"9D",x"00",x"CD",x"B2",x"27",x"27",x"49",x"B1",x"AA",x"2C",x"D2",x"8C",x"EC",x"31",x"BC",x"27",x"EE",x"30",x"92",x"B1",x"B0",x"E8",x"2A",x"C3",x"8A",x"B2",x"43",x"A5",x"26",x"0F",x"3B",x"B1",x"2E",x"23",x"BF",x"3D",x"EC",x"C4",x"BA",x"8C",x"FC",x"CE",x"70",x"12",x"ED",x"32",x"B2",x"B9",x"CD",x"4D",x"B8",x"DB",x"44",x"E6",x"36",x"3F",x"A8",x"4A",x"53",x"B3",x"5F",x"92",x"24",x"52",x"23",x"7C",x"4A",x"B0",x"92",x"C8",x"70",x"CE",x"C9",x"CE",x"4A",x"AC",x"2A",x"C8",x"6F",x"1B",x"3B",x"B1",x"4D",x"92",x"78",x"EA",x"9C",x"48",x"BB",x"8C",x"6D",x"2E",x"0A",x"6A",x"30",x"96",x"A8",x"31",x"C3",x"AF",x"49",x"C4",x"B2",x"AA",x"0E",x"37",x"07",x"8E",x"98",x"8E",x"33",x"BC",x"52",x"38",x"74",x"CA",x"F1",x"88",x"72",x"E1",x"8A",x"0D",x"C7",x"2D",x"2A",x"59",x"53",x"B7",x"E5",x"A4",x"A0",x"14",x"33",x"CB",x"B6",x"4A",x"80",x"64",x"54",x"8D",x"5F",x"A3",x"8A",x"44",x"55",x"35",x"6E",x"8E",x"EC",x"31",x"15",x"DB",x"78",x"A5",x"88",x"5B",x"B7",x"63",x"02",x"84",x"C2",x"43",x"80",x"98",x"A5",x"31",x"F0",x"00",x"FF",
		x"60",x"A1",x"88",x"9D",x"D2",x"C8",x"BB",x"8C",x"B8",x"0C",x"0E",x"76",x"ED",x"3C",x"C2",x"96",x"4C",x"29",x"7D",x"F1",x"08",x"6B",x"51",x"15",x"F7",x"96",x"21",x"A8",x"9E",x"A4",x"29",x"6B",x"B7",x"A0",x"06",x"53",x"37",x"6D",x"34",x"82",x"92",x"5C",x"D5",x"73",x"F1",x"08",x"4B",x"72",x"33",x"AB",x"BA",x"23",x"2A",x"31",x"D5",x"2D",x"E7",x"8C",x"38",x"A7",x"30",x"53",x"6D",x"D2",x"E2",x"1A",x"55",x"43",x"24",x"55",x"4A",x"4A",x"60",x"69",x"92",x"CC",x"2C",x"4F",x"8E",x"B9",x"D9",x"D2",x"8E",x"B2",x"24",x"55",x"0B",x"8B",x"3B",x"CA",x"5C",x"45",x"3D",x"B9",x"DD",x"A8",x"73",x"77",x"B1",x"E0",x"B4",x"AD",x"CE",x"53",x"34",x"9C",x"DA",x"B4",x"3A",x"4F",x"B6",x"74",x"5E",x"5D",x"9A",x"34",x"D0",x"CB",x"74",x"55",x"6A",x"F3",x"C1",x"0C",x"D1",x"45",x"66",x"CA",x"15",x"3D",x"DC",x"1B",x"A9",x"22",x"35",x"51",x"4F",x"DA",x"62",x"AA",x"DC",x"55",x"3C",x"B9",x"B7",x"AA",x"F3",x"14",x"4D",x"A3",x"CE",x"AA",x"CE",x"53",x"34",x"9D",x"BB",x"A8",x"26",x"0D",x"B2",x"52",x"6B",x"03",x"00",x"90",x"A2",x"A6",x"44",x"3D",x"7C",x"61",x"F3",x"53",x"A6",x"B4",x"EA",x"A8",x"CD",x"8D",x"C9",x"D3",x"2C",x"C6",x"36",x"27",x"D4",x"0A",x"76",x"AF",x"DD",x"2C",x"9F",x"26",x"D9",x"25",x"71",x"31",x"74",x"E9",x"54",x"53",x"25",x"41",x"53",x"39",x"4B",x"24",x"ED",x"08",x"2B",x"0A",x"0D",x"53",x"0B",x"A3",x"FC",x"94",x"D9",x"AD",x"2A",x"8A",x"F2",x"62",x"F6",x"30",x"CF",x"B1",x"CE",x"29",x"DC",x"3B",x"DD",x"E4",x"28",x"60",x"7B",x"11",x"03",x"AC",x"56",x"AA",x"80",x"35",x"DB",x"14",x"30",x"EB",x"94",x"00",x"C6",x"CC",x"2C",x"4E",x"CD",x"C2",x"A2",x"3E",x"A7",x"B8",x"59",x"B8",x"6A",x"C9",x"92",x"E2",x"26",x"AE",x"E1",x"2E",x"4D",x"93",x"5B",x"B9",x"58",x"98",x"C6",x"05",x"01",x"34",x"E7",x"C1",x"80",x"16",x"D5",x"09",x"E0",x"35",x"3B",x"01",x"84",x"D5",x"40",x"40",x"94",x"6E",x"08",x"28",x"CE",x"94",x"01",x"25",x"85",x"3B",x"AF",x"58",x"F7",x"14",x"71",x"52",x"C2",x"98",x"2D",x"85",x"74",x"69",x"09",x"63",x"B4",x"30",x"D6",x"A5",x"25",x"0E",x"DE",x"DC",x"C5",x"96",x"86",x"D4",x"67",x"53",x"93",x"78",x"52",x"0A",x"1B",x"2C",x"5C",x"63",x"4D",x"A9",x"BC",x"B1",x"68",x"D5",x"B6",x"A5",x"F5",x"26",x"3C",x"C5",x"BA",x"A6",x"DE",x"DB",x"88",x"10",x"CB",x"9A",x"A6",x"68",x"35",x"83",x"A4",x"6B",x"58",x"A2",x"0B",x"37",x"96",x"A4",x"66",x"89",x"C9",x"52",x"49",x"3B",x"B3",x"3C",x"58",x"C9",x"14",x"DD",x"22",x"AA",x"18",x"D9",x"5C",x"BD",x"2D",x"AA",x"BD",x"0A",x"2B",x"B3",x"B4",x"62",x"AB",x"5E",x"9C",x"65",x"62",x"D1",x"ED",x"01",x"FF",
		x"60",x"0C",x"38",x"22",x"43",x"00",x"4B",x"A5",x"09",x"60",x"AB",x"F6",x"96",x"0E",x"95",x"62",x"62",x"8D",x"5B",x"94",x"13",x"B9",x"CF",x"C4",x"1D",x"71",x"4B",x"2A",x"EA",x"53",x"77",x"84",x"D5",x"91",x"79",x"6D",x"9D",x"11",x"B4",x"28",x"14",x"D9",x"55",x"46",x"D0",x"1C",x"53",x"55",x"45",x"19",x"61",x"35",x"4C",x"D3",x"19",x"75",x"84",x"55",x"93",x"54",x"4F",x"98",x"11",x"B6",x"C0",x"1C",x"DE",x"55",x"5A",x"D2",x"BC",x"B1",x"79",x"55",x"49",x"51",x"F3",x"22",x"96",x"5D",x"27",x"04",x"2D",x"08",x"5B",x"66",x"12",x"17",x"34",x"4F",x"1C",x"39",x"61",x"42",x"D8",x"9D",x"9A",x"BA",x"39",x"35",x"E1",x"50",x"22",x"5A",x"19",x"87",x"00",x"2B",x"99",x"08",x"60",x"48",x"B6",x"64",x"57",x"41",x"92",x"ED",x"B6",x"87",x"DD",x"1D",x"63",x"4D",x"5A",x"6E",x"F6",x"10",x"82",x"B9",x"69",x"A6",x"B9",x"5D",x"09",x"F6",x"86",x"95",x"E6",x"75",x"43",x"58",x"95",x"76",x"46",x"30",x"9D",x"A1",x"75",x"C5",x"6E",x"F1",x"D4",x"82",x"3E",x"6D",x"A7",x"A5",x"43",x"0A",x"C6",x"76",x"DC",x"91",x"0F",x"23",x"E8",x"3D",x"71",x"46",x"35",x"8C",x"A0",x"75",x"C7",x"1E",x"75",x"B7",x"8A",x"16",x"5B",x"7B",x"B4",x"DD",x"19",x"9A",x"DE",x"9C",x"D6",x"0F",x"57",x"68",x"30",x"B3",x"5D",x"38",x"A4",x"91",x"6B",x"A4",x"72",x"E9",x"52",x"CD",x"C2",x"DA",x"C8",x"E5",x"4B",x"07",x"99",x"68",x"6A",x"57",x"4C",x"5D",x"A2",x"AC",x"89",x"5C",x"3D",x"4C",x"90",x"91",x"A7",x"26",x"40",x"0F",x"8A",x"04",x"08",x"5C",x"05",x"18",x"D0",x"B5",x"5B",x"4A",x"4B",x"30",x"36",x"B1",x"B4",x"2D",x"0F",x"51",x"52",x"B8",x"DB",x"B4",x"DC",x"FB",x"32",x"67",x"DB",x"52",x"AA",x"C8",x"27",x"53",x"29",x"77",x"E9",x"82",x"BA",x"72",x"A6",x"DE",x"AD",x"C9",x"64",x"BA",x"1C",x"72",x"8F",x"32",x"CA",x"2B",x"13",x"EA",x"3C",x"F2",x"A0",x"AE",x"54",x"B8",x"F3",x"C8",x"82",x"BA",x"16",x"E1",x"CC",x"2D",x"F3",x"6A",x"DB",x"44",x"52",x"99",x"3A",x"B0",x"8E",x"50",x"4E",x"4D",x"80",x"A0",x"2E",x"47",x"5C",x"5D",x"A4",x"9A",x"39",x"1D",x"69",x"0E",x"1E",x"62",x"51",x"67",x"E4",x"29",x"9A",x"B1",x"67",x"ED",x"91",x"27",x"6D",x"19",x"EA",x"66",x"5A",x"9E",x"B4",x"84",x"79",x"DA",x"2E",x"65",x"52",x"1C",x"66",x"65",x"27",x"D4",x"5E",x"72",x"A7",x"66",x"94",x"50",x"5B",x"69",x"61",x"91",x"89",x"A1",x"95",x"C3",x"A7",x"49",x"48",x"9C",x"51",x"A4",x"2C",x"26",x"56",x"75",x"46",x"19",x"B2",x"85",x"AA",x"2D",x"1E",x"A5",x"4B",x"ED",x"AA",x"D6",x"B9",x"55",x"B6",x"8C",x"AB",x"58",x"D7",x"51",x"DB",x"32",x"66",x"22",x"5D",x"46",x"EB",x"43",x"45",x"0B",x"76",x"1E",x"9D",x"8F",x"65",x"15",x"D4",x"75",x"8C",x"D1",x"97",x"64",x"63",x"EE",x"31",x"A7",x"18",x"D2",x"8D",x"9D",x"DB",x"9A",x"AA",x"4A",x"17",x"2E",x"69",x"6B",x"AA",x"A2",x"9D",x"B4",x"A6",x"AC",x"A9",x"92",x"75",x"C8",x"E6",x"B6",x"E4",x"62",x"1C",x"A1",x"AB",x"DB",x"56",x"6C",x"18",x"6B",x"4C",x"2E",x"7B",x"36",x"61",x"6E",x"55",x"36",x"ED",x"C9",x"86",x"7A",x"46",x"B8",x"B0",x"67",x"5F",x"EC",x"2D",x"CE",x"08",x"10",x"62",x"30",x"03",x"A2",x"0F",x"26",x"40",x"54",x"25",x"04",x"48",x"BC",x"19",x"01",x"5E",x"95",x"3E",x"FF",
		x"60",x"04",x"18",x"24",x"9D",x"01",x"5B",x"8D",x"09",x"60",x"E8",x"D1",x"12",x"E6",x"C4",x"EA",x"B9",x"71",x"5B",x"98",x"23",x"8B",x"E7",x"D6",x"1D",x"41",x"8D",x"C2",x"51",x"5B",x"65",x"04",x"3D",x"2A",x"AB",x"4D",x"ED",x"11",x"F4",x"C4",x"AC",x"D1",x"75",x"5A",x"D8",x"82",x"8B",x"7A",x"C4",x"2E",x"61",x"B3",x"AD",x"6A",x"62",x"2B",x"85",x"D5",x"BB",x"5A",x"44",x"9C",x"10",x"B4",x"A0",x"62",x"5E",x"71",x"5D",x"D0",x"A3",x"88",x"5A",x"C7",x"B1",x"01",x"03",x"9A",x"57",x"2F",x"7E",x"88",x"95",x"61",x"52",x"B5",x"78",x"3E",x"75",x"AA",x"D8",x"ED",x"E2",x"85",x"54",x"29",x"6C",x"57",x"8A",x"17",x"82",x"17",x"B3",x"4F",x"09",x"41",x"CA",x"A2",x"E2",x"11",x"87",x"01",x"7D",x"4D",x"0B",x"60",x"F4",x"49",x"01",x"8C",x"DA",x"95",x"B2",x"6E",x"D5",x"32",x"23",x"52",x"29",x"4A",x"E0",x"A0",x"4D",x"AB",x"A5",x"4C",x"4E",x"42",x"A3",x"C4",x"96",x"3A",x"59",x"0E",x"8E",x"72",x"52",x"9A",x"62",x"D9",x"D9",x"DD",x"4D",x"6A",x"AB",x"25",x"13",x"33",x"37",x"A9",x"AB",x"9A",x"4C",x"D5",x"93",x"84",x"AE",x"48",x"32",x"D7",x"AC",x"8D",x"80",x"25",x"DD",x"05",x"50",x"61",x"AA",x"00",x"B6",x"AE",x"54",x"40",x"31",x"2A",x"04",x"28",x"5A",x"94",x"01",x"5A",x"AB",x"A7",x"34",x"5A",x"4F",x"77",x"B3",x"9D",x"32",x"3B",x"C2",x"83",x"A5",x"4D",x"C9",x"5D",x"2D",x"2D",x"A3",x"CC",x"25",x"F7",x"CD",x"6C",x"94",x"BB",x"94",x"3C",x"54",x"F1",x"16",x"6D",x"53",x"8A",x"98",x"D9",x"9B",x"7D",x"49",x"2A",x"82",x"4E",x"57",x"8D",x"3A",x"A9",x"48",x"D4",x"23",x"C8",x"67",x"8F",x"B4",x"F8",x"54",x"91",x"A9",x"32",x"E2",x"E2",x"45",x"3C",x"37",x"EC",x"88",x"5A",x"64",x"B1",x"98",x"38",x"23",x"6C",x"89",x"45",x"63",x"A3",x"A0",x"30",x"7B",x"E7",x"94",x"B0",x"3A",x"A2",x"16",x"C5",x"28",x"B3",x"CE",x"08",x"6B",x"67",x"D5",x"F0",x"D9",x"2D",x"2A",x"93",x"34",x"CC",x"16",x"97",x"A4",x"0C",x"34",x"D3",x"58",x"9A",x"D2",x"36",x"88",x"CD",x"B3",x"4E",x"AA",x"5A",x"62",x"D1",x"98",x"38",x"26",x"AB",x"86",x"D8",x"AB",x"E2",x"94",x"A4",x"57",x"25",x"D1",x"AC",x"DB",x"C2",x"96",x"19",x"CD",x"73",x"4E",x"0B",x"6B",x"64",x"51",x"CB",x"39",x"2D",x"CA",x"9E",x"5D",x"B4",x"A6",x"94",x"24",x"1A",x"49",x"B1",x"9C",x"13",x"2A",x"6F",x"35",x"D9",x"AB",x"96",x"E9",x"9C",x"D1",x"72",x"EB",x"46",x"62",x"2A",x"5E",x"55",x"D4",x"EB",x"22",x"60",x"84",x"46",x"15",x"76",x"ED",x"68",x"EE",x"AB",x"4C",x"34",x"58",x"B2",x"99",x"67",x"51",x"C9",x"E0",x"21",x"26",x"9A",x"84",x"00",x"81",x"96",x"11",x"A0",x"C0",x"50",x"04",x"34",x"E2",x"F6",x"00",x"FF",
		x"60",x"04",x"E8",x"2A",x"43",x"00",x"CB",x"64",x"08",x"60",x"29",x"8F",x"14",x"84",x"2C",x"11",x"A2",x"9D",x"52",x"68",x"BA",x"65",x"89",x"2C",x"49",x"81",x"ED",x"EE",x"AD",x"D4",x"AE",x"F8",x"BE",x"B9",x"B6",x"73",x"BA",x"E2",x"C7",x"AA",x"96",x"A9",x"E9",x"4A",x"98",x"0B",x"5B",x"B9",x"35",x"11",x"C0",x"C8",x"E9",x"0C",x"B8",x"D1",x"5C",x"00",x"93",x"72",x"09",x"60",x"72",x"CE",x"36",x"65",x"6B",x"1E",x"EE",x"4D",x"D2",x"94",x"06",x"66",x"68",x"2C",x"2E",x"6D",x"AC",x"98",x"A9",x"9A",x"BA",x"B5",x"A1",x"B2",x"47",x"78",x"B2",x"D2",x"C6",x"26",x"52",x"49",x"5D",x"4B",x"17",x"9B",x"48",x"15",x"75",x"29",x"5D",x"EA",x"22",x"D1",x"D4",x"A5",x"F4",x"69",x"B2",x"56",x"70",x"97",x"D2",x"E5",x"89",x"EE",x"AE",x"AB",x"5A",x"97",x"12",x"B9",x"67",x"64",x"6A",x"5D",x"31",x"16",x"6C",x"DE",x"48",x"00",x"5B",x"45",x"0A",x"60",x"B0",x"8C",x"D0",x"C4",x"CA",x"E2",x"21",x"89",x"43",x"91",x"0A",x"B9",x"48",x"C7",x"1D",x"69",x"C9",x"AA",x"6A",x"39",x"67",x"A4",x"35",x"AA",x"58",x"74",x"ED",x"91",x"B6",x"C0",x"62",x"35",x"71",x"46",x"DA",x"04",x"6B",x"56",x"57",x"19",x"59",x"B3",x"4C",x"56",x"35",x"4A",x"E4",x"5E",x"9A",x"67",x"A8",x"6D",x"54",x"05",x"A9",x"56",x"A1",x"89",x"46",x"32",x"9A",x"0A",x"49",x"24",x"1D",x"D1",x"34",x"46",x"A2",x"9D",x"74",x"84",x"D3",x"18",x"B2",x"6F",x"92",x"12",x"36",x"2E",x"94",x"D3",x"4E",x"4A",x"50",x"85",x"50",x"CF",x"D8",x"0A",x"49",x"37",x"44",x"B6",x"EB",x"C4",x"B5",x"45",x"A2",x"D5",x"A4",x"9D",x"52",x"36",x"4D",x"EA",x"3D",x"49",x"5B",x"D0",x"03",x"8B",x"E6",x"54",x"1E",x"41",x"73",x"A2",x"12",x"53",x"A5",x"84",x"49",x"A9",x"45",x"94",x"AD",x"12",x"15",x"49",x"65",x"DE",x"0C",x"43",x"14",x"94",x"94",x"5B",x"D1",x"32",x"49",x"50",x"EA",x"1E",x"91",x"50",x"15",x"89",x"93",x"67",x"7A",x"92",x"54",x"B7",x"20",x"AE",x"6A",x"4E",x"47",x"54",x"12",x"2B",x"FB",x"24",x"1E",x"61",x"CD",x"A2",x"1C",x"53",x"65",x"F8",x"35",x"A8",x"B2",x"6E",x"9C",x"E9",x"B7",x"68",x"C9",x"75",x"11",x"4B",x"2C",x"80",x"49",x"9D",x"5B",x"BC",x"45",x"88",x"99",x"C5",x"1E",x"71",x"F2",x"EA",x"E2",x"1B",x"77",x"14",x"C9",x"B9",x"9B",x"5A",x"9D",x"52",x"16",x"27",x"2A",x"3E",x"51",x"58",x"55",x"AA",x"0A",x"C6",x"DA",x"19",x"5D",x"62",x"DD",x"26",x"BC",x"78",x"0C",x"89",x"75",x"9B",x"C8",x"92",x"36",x"26",x"3E",x"AD",x"6C",x"73",x"DB",x"1C",x"E5",x"BA",x"A5",x"95",x"2B",x"4B",x"62",x"E3",x"16",x"36",x"39",x"AC",x"C1",x"BC",x"52",x"44",x"55",x"B5",x"F9",x"F8",x"C2",x"56",x"55",x"D5",x"16",x"E5",x"B5",x"92",x"37",x"55",x"7B",x"C6",x"D3",x"4E",x"B2",x"98",x"1D",x"51",x"4C",x"AB",x"D8",x"DC",x"07",x"FF",
		x"60",x"08",x"68",x"55",x"9D",x"01",x"63",x"8D",x"0B",x"60",x"F4",x"29",x"03",x"F4",x"19",x"D1",x"BC",x"52",x"C4",x"CD",x"BD",x"4E",x"0B",x"52",x"AA",x"08",x"8D",x"39",x"CD",x"8F",x"65",x"CC",x"32",x"6B",x"37",x"3F",x"95",x"74",x"8B",x"AA",x"D3",x"FC",x"5C",x"3C",x"CC",x"BB",x"6E",x"0B",x"4B",x"B0",x"A4",x"EC",x"A6",x"02",x"A8",x"06",x"45",x"79",x"35",x"A9",x"AA",x"5B",x"9D",x"14",x"14",x"3D",x"1E",x"1A",x"69",x"53",x"30",x"58",x"55",x"86",x"25",x"0D",x"7E",x"15",x"DB",x"AA",x"B1",x"D4",x"F8",x"B9",x"7A",x"68",x"74",x"1D",x"04",x"84",x"A4",x"99",x"BC",x"59",x"DC",x"D5",x"D4",x"72",x"09",x"4A",x"21",x"63",x"B7",x"CD",x"2D",x"C8",x"91",x"5C",x"5D",x"BA",x"94",x"30",x"17",x"72",x"13",x"77",x"57",x"82",x"92",x"25",x"18",x"AB",x"76",x"F3",x"73",x"90",x"D4",x"C8",x"3A",x"C3",x"CB",x"29",x"5C",x"3D",x"AB",x"0C",x"27",x"15",x"0F",x"F5",x"AA",x"DA",x"AC",x"D4",x"2C",x"2C",x"BA",x"6C",x"B3",x"72",x"D2",x"92",x"EC",x"A8",x"C6",x"2E",x"51",x"42",x"A2",x"22",x"97",x"A0",x"BB",x"70",x"56",x"8F",x"5C",x"82",x"9A",x"D4",x"C4",x"AD",x"49",x"F1",x"4A",x"35",x"37",x"F7",x"3A",x"CD",x"CD",x"D9",x"CC",x"D2",x"C2",x"34",x"37",x"37",x"D6",x"4C",x"A9",x"5A",x"DC",x"DC",x"29",x"DC",x"B4",x"59",x"71",x"F3",x"C0",x"32",x"8E",x"36",x"C9",x"CD",x"07",x"DD",x"CD",x"D2",x"30",x"A0",x"15",x"09",x"06",x"D4",x"AC",x"56",x"B2",x"12",x"C4",x"BC",x"AB",x"CE",x"C8",x"4A",x"63",x"F3",x"9C",x"38",x"23",x"2D",x"55",x"DC",x"AA",x"AD",x"B6",x"38",x"46",x"B3",x"8C",x"B2",x"EA",x"F2",x"DC",x"51",x"23",x"D2",x"59",x"8B",x"B2",x"77",x"35",x"E9",x"38",x"2B",x"4E",x"51",x"DC",x"A2",x"16",x"B7",x"34",x"0F",x"4A",x"63",x"5F",x"55",x"B2",x"D8",x"29",x"5C",x"2D",x"6D",x"A8",x"4A",x"15",x"B7",x"EC",x"38",x"C0",x"80",x"E2",x"24",x"08",x"90",x"24",x"54",x"8A",x"8A",x"72",x"57",x"8F",x"36",x"25",x"8C",x"DE",x"CD",x"D3",x"6C",x"8F",x"20",x"86",x"34",x"CB",x"88",x"32",x"C2",x"98",x"4A",x"35",x"AB",x"CA",x"08",x"4B",x"70",x"53",x"CF",x"D9",x"23",x"AC",x"C9",x"54",x"3D",x"E7",x"8C",x"A8",x"46",x"65",x"CF",x"9A",x"33",x"B2",x"5A",x"8D",x"D5",x"63",x"F5",x"A8",x"6A",x"74",x"D2",x"F2",x"4E",x"AD",x"2B",x"D9",x"C9",x"4A",x"7A",x"B7",x"A1",x"14",x"23",x"6B",x"EE",x"5D",x"C6",x"DC",x"95",x"B5",x"A4",x"6D",x"99",x"4A",x"57",x"91",x"D4",x"B6",x"69",x"A9",x"C1",x"58",x"2B",x"3A",x"A7",x"A5",x"85",x"16",x"4E",x"F7",x"5A",x"96",x"E6",x"5A",x"38",x"BC",x"19",x"01",x"A2",x"77",x"22",x"40",x"4C",x"A4",x"04",x"88",x"11",x"03",x"01",x"2E",x"70",x"20",x"80",x"85",x"08",x"00",x"00",x"80",x"30",x"4D",x"AD",x"82",x"56",x"8D",x"DB",x"30",x"BD",x"29",x"72",x"2E",x"19",x"6D",x"F7",x"21",x"A8",x"B9",x"66",x"D4",x"2D",x"86",x"88",x"D5",x"92",x"51",x"55",x"9F",x"62",x"51",x"4B",x"46",x"5D",x"6D",x"AA",x"47",x"2E",x"19",x"7D",x"09",x"C5",x"16",x"35",x"07",x"08",x"10",x"84",x"07",x"03",x"A2",x"14",x"33",x"75",x"F3",x"21",x"62",x"B9",x"C4",x"55",x"CD",x"96",x"A8",x"57",x"13",x"D7",x"34",x"DD",x"62",x"11",x"4B",x"54",x"5B",x"5D",x"89",x"79",x"4F",x"25",x"80",x"0F",x"E6",x"0F",x"FF",
		x"60",x"08",x"28",x"3E",x"8C",x"00",x"C5",x"BA",x"13",x"A0",x"58",x"37",x"D7",x"FA",x"95",x"2E",x"3A",x"71",x"52",x"17",x"46",x"87",x"C8",x"CC",x"2E",x"43",x"A8",x"E3",x"EA",x"55",x"BB",x"0C",x"B1",x"8C",x"69",x"56",x"ED",x"D6",x"67",x"5F",x"AD",x"16",x"75",x"5A",x"D7",x"7C",x"8C",x"99",x"37",x"69",x"6D",x"0F",x"99",x"EC",x"36",x"A7",x"35",x"3D",x"A4",x"52",x"C4",x"E4",x"56",x"77",x"E9",x"2C",x"95",x"41",x"4A",x"95",x"71",x"B9",x"26",x"3B",x"29",x"65",x"22",x"ED",x"EA",x"EA",x"B8",x"55",x"99",x"96",x"99",x"6A",x"E2",x"56",x"15",x"A5",x"2E",x"6C",x"71",x"5A",x"D5",x"AC",x"3A",x"A9",x"56",x"2E",x"6D",x"F7",x"A1",x"E8",x"3E",x"B9",x"35",x"DD",x"A9",x"B0",x"66",x"95",x"96",x"75",x"A3",x"4C",x"59",x"93",x"5B",x"D6",x"AD",x"31",x"46",x"4F",x"6E",x"D9",x"34",x"22",x"E4",x"35",x"AB",x"E5",x"C3",x"29",x"63",x"F6",x"E4",x"96",x"37",x"27",x"24",x"57",x"B3",x"5B",x"51",x"BD",x"88",x"75",x"35",x"1A",x"65",x"8D",x"2A",x"11",x"D3",x"78",x"14",x"35",x"86",x"A4",x"D7",x"9C",x"96",x"97",x"A4",x"D2",x"D1",x"53",x"42",x"5E",x"83",x"51",x"44",x"2C",x"76",x"79",x"F7",x"21",x"68",x"DE",x"34",x"E5",x"D5",x"A9",x"68",x"69",x"D2",x"51",x"54",x"3F",x"EE",x"2A",x"4E",x"46",x"39",x"4C",x"A8",x"46",x"35",x"1E",x"45",x"37",x"25",x"16",x"D9",x"86",x"01",x"4D",x"37",x"97",x"7C",x"A8",x"E2",x"D0",x"9C",x"5D",x"FA",x"64",x"25",x"BC",x"36",x"D4",x"98",x"53",x"50",x"9E",x"EA",x"A8",x"65",x"C9",x"5E",x"42",x"73",x"ED",x"B8",x"2B",x"2B",x"57",x"CF",x"A9",x"0C",x"08",x"68",x"3A",x"0C",x"01",x"15",x"76",x"22",x"20",x"A1",x"75",x"04",x"78",x"EB",x"89",x"00",x"6F",x"3D",x"1E",x"FF",
		x"60",x"08",x"A8",x"D5",x"BC",x"14",x"35",x"BA",x"87",x"7B",x"E9",x"16",x"E7",x"62",x"EE",x"D1",x"55",x"5B",x"54",x"A2",x"4B",x"C4",x"4C",x"6D",x"71",x"B5",x"2E",x"EE",x"35",x"A5",x"E4",x"4D",x"06",x"9B",x"C6",x"E4",x"52",x"2D",x"97",x"AA",x"82",x"4E",x"5A",x"D2",x"62",x"8A",x"A2",x"57",x"6E",x"5E",x"8F",x"46",x"2C",x"3D",x"B7",x"D9",x"D3",x"38",x"89",x"65",x"94",x"66",x"76",x"EE",x"6C",x"E1",x"51",x"92",x"31",x"94",x"91",x"99",x"A7",x"01",x"04",x"30",x"5E",x"E9",x"C2",x"C4",x"8D",x"D3",x"2B",x"52",x"09",x"B2",x"62",x"CB",x"28",x"B3",x"2D",x"2A",x"52",x"BC",x"2D",x"22",x"B7",x"38",x"29",x"F1",x"D2",x"8C",x"D3",x"E2",x"6C",x"C5",x"43",x"2B",x"76",x"CB",x"92",x"C9",x"0C",x"F1",x"56",x"25",x"4D",x"FA",x"DA",x"45",x"3B",x"95",x"24",x"EA",x"6B",x"13",x"6B",x"5D",x"A2",x"E0",x"AE",x"5C",x"AC",x"69",x"09",x"7D",x"F8",x"30",x"C9",x"BA",x"29",x"0E",x"EE",x"DC",x"29",x"E3",x"A4",x"34",x"AB",x"B6",x"14",x"AF",x"55",x"A2",x"2C",x"3B",x"42",x"DC",x"76",x"89",x"A2",x"EA",x"70",x"F1",x"D9",x"29",x"8E",x"AA",x"D3",x"59",x"6F",x"97",x"38",x"9A",x"AD",x"30",x"8B",x"13",x"A2",x"68",x"3B",x"2A",x"C3",x"36",x"02",x"8A",x"72",x"47",x"40",x"F1",x"A1",x"04",x"C8",x"CE",x"D5",x"38",x"26",x"BB",x"99",x"55",x"AD",x"64",x"3A",x"EF",x"69",x"E2",x"B5",x"93",x"E5",x"BC",x"A7",x"89",x"CF",x"0E",x"AE",x"F1",x"11",x"2E",x"BE",x"38",x"F8",x"C6",x"97",x"9B",x"DA",x"A2",x"10",x"9B",x"E8",x"A1",x"92",x"B5",x"43",x"E6",x"A3",x"AA",x"49",x"36",x"0E",x"75",x"8A",x"AA",x"26",x"DE",x"18",x"D5",x"99",x"9B",x"3A",x"7B",x"ED",x"D6",x"6D",x"14",x"2E",x"46",x"AD",x"DA",x"70",x"60",x"26",x"2B",x"ED",x"6E",x"C3",x"60",x"19",x"29",x"BC",x"A4",x"8D",x"5D",x"97",x"3B",x"D9",x"D2",x"36",x"B5",x"D0",x"22",x"94",x"4B",x"DA",x"34",x"62",x"A9",x"60",x"AC",x"69",x"F3",x"48",x"29",x"42",x"D1",x"1A",x"08",x"90",x"50",x"59",x"E8",x"06",x"A9",x"70",x"C1",x"25",x"6D",x"EC",x"3C",x"CD",x"59",x"67",x"B7",x"A9",x"CB",x"52",x"13",x"9B",x"DA",x"96",x"6E",x"53",x"9D",x"7D",x"59",x"5B",x"9B",x"33",x"51",x"E9",x"35",x"6D",x"6D",x"DE",x"98",x"AD",x"57",x"97",x"AD",x"6B",x"56",x"C9",x"9A",x"95",x"F6",x"EE",x"55",x"D0",x"AB",x"8E",x"BD",x"1E",x"FF",
		x"60",x"2D",x"18",x"3E",x"4D",x"54",x"D4",x"8C",x"A8",x"1A",x"4D",x"4D",x"DF",x"32",x"C2",x"62",x"3D",x"A5",x"62",x"CD",x"F0",x"9B",x"B7",x"54",x"B7",x"C5",x"C3",x"AF",x"CE",x"82",x"DD",x"EE",x"04",x"BF",x"44",x"0B",x"B6",x"C8",x"D2",x"82",x"98",x"38",x"33",x"BD",x"4D",x"0B",x"63",x"61",x"F7",x"B2",x"74",x"2D",x"4E",x"CD",x"D4",x"CD",x"9C",x"B5",x"38",x"9A",x"E6",x"70",x"6D",x"D6",x"E2",x"24",x"DA",x"C2",x"65",x"EE",x"88",x"B2",x"CE",x"70",x"F1",x"6A",x"23",x"4A",x"6E",x"DC",x"2C",x"EE",x"8C",x"38",x"9B",x"71",x"37",x"BF",x"33",x"92",x"2A",x"DB",x"53",x"ED",x"71",x"C8",x"6B",x"8A",x"50",x"B6",x"2C",x"08",x"D0",x"B1",x"4D",x"45",x"C9",x"4E",x"98",x"C5",x"63",x"13",x"27",x"37",x"E1",x"9C",x"77",x"4C",x"52",x"65",x"47",x"AA",x"DD",x"16",x"B9",x"57",x"52",x"6B",x"52",x"C7",x"94",x"D9",x"88",x"BA",x"44",x"6B",x"57",x"24",x"45",x"3E",x"AE",x"65",x"4B",x"DE",x"55",x"88",x"1A",x"3F",x"1A",x"79",x"B3",x"61",x"66",x"FE",x"78",x"94",x"D5",x"A7",x"4B",x"C4",x"92",x"56",x"D7",x"64",x"2E",x"61",x"6B",x"52",x"D3",x"56",x"2A",x"BB",x"E4",x"06",x"02",x"94",x"C9",x"4E",x"80",x"29",x"47",x"10",x"B0",x"55",x"31",x"02",x"26",x"77",x"01",x"02",x"4C",x"E6",x"56",x"FA",x"EC",x"BC",x"39",x"63",x"4A",x"1B",x"AA",x"B5",x"51",x"B7",x"CD",x"6D",x"AC",x"D6",x"46",x"DD",x"37",x"F7",x"A9",x"4D",x"D5",x"DA",x"A8",x"7B",x"97",x"B6",x"54",x"E7",x"C3",x"11",x"9B",x"DB",x"D2",x"BC",x"8F",x"BA",x"6E",x"6E",x"6B",x"8F",x"31",x"6A",x"BC",x"B8",x"6D",x"35",x"66",x"72",x"D8",x"94",x"B6",x"57",x"17",x"C9",x"E9",x"93",x"CB",x"5E",x"AD",x"B7",x"B8",x"36",x"2A",x"47",x"73",x"D6",x"6C",x"DA",x"B0",x"9E",x"E9",x"2A",x"CE",x"92",x"C3",x"2A",x"BA",x"3B",x"39",x"0D",x"49",x"0F",x"29",x"EF",x"07",x"FF",
		x"60",x"A1",x"AE",x"46",x"5C",x"3D",x"BB",x"94",x"7A",x"14",x"4D",x"76",x"DA",x"32",x"AA",x"91",x"AD",x"C8",x"79",x"F5",x"28",x"7B",x"D2",x"22",x"D3",x"D5",x"A3",x"68",x"41",x"13",x"23",x"56",x"9B",x"A2",x"59",x"4E",x"F6",x"58",x"33",x"F2",x"61",x"25",x"C4",x"65",x"ED",x"C8",x"AB",x"37",x"E7",x"D0",x"AD",x"23",x"2B",x"C9",x"8D",x"8A",x"DB",x"B5",x"B4",x"D4",x"50",x"6A",x"4E",x"DB",x"E2",x"D2",x"4D",x"64",x"A8",x"5B",x"4B",x"73",x"17",x"D5",x"96",x"B6",x"A5",x"C8",x"9D",x"DC",x"DA",x"9A",x"96",x"2A",x"77",x"11",x"69",x"69",x"53",x"AA",x"32",x"4C",x"B5",x"29",x"61",x"29",x"F2",x"22",x"8D",x"94",x"D6",x"25",x"CD",x"93",x"2C",x"93",x"16",x"97",x"38",x"8F",x"60",x"69",x"F2",x"56",x"82",x"DC",x"9C",x"75",x"29",x"6B",x"F1",x"73",x"0B",x"96",x"65",x"AF",x"C9",x"4F",x"CB",x"D5",x"1A",x"BD",x"96",x"20",x"2D",x"53",x"6F",x"48",x"5B",x"C2",x"D4",x"55",x"A2",x"39",x"6B",x"89",x"F3",x"60",x"F1",x"92",x"2D",x"25",x"2D",x"C1",x"99",x"CB",x"BB",x"B4",x"AC",x"2A",x"71",x"89",x"AC",x"D3",x"B2",x"A6",x"D5",x"28",x"B2",x"4E",x"CB",x"9B",x"73",x"45",x"AF",x"26",x"A5",x"E8",x"DE",x"14",x"35",x"1B",x"A7",x"B2",x"1B",x"31",x"CA",x"5C",x"AC",x"AA",x"6E",x"4C",x"C9",x"BB",x"C9",x"03",x"FF",
		x"60",x"04",x"98",x"A4",x"8C",x"00",x"DD",x"66",x"94",x"A4",x"A6",x"4A",x"D7",x"AC",x"DD",x"C2",x"E2",x"3A",x"DD",x"A2",x"F6",x"F0",x"8B",x"DC",x"74",x"F7",x"D9",x"C3",x"29",x"EA",x"42",x"23",x"EA",x"0C",x"3B",x"87",x"35",x"CB",x"88",x"33",x"EC",x"12",x"DB",x"DD",x"33",x"CA",x"70",x"6B",x"CC",x"74",x"C9",x"32",x"C3",x"AD",x"A5",x"DD",x"39",x"AA",x"0C",x"B7",x"8D",x"74",x"96",x"A8",x"33",x"BC",x"9E",x"92",x"55",x"B2",x"CA",x"F0",x"87",x"0F",x"72",x"CB",x"32",x"C5",x"1F",x"C6",x"D1",x"A2",x"66",x"15",x"BF",x"18",x"91",x"B6",x"48",x"92",x"FC",x"EA",x"48",x"8B",x"32",x"4E",x"0A",x"B3",x"61",x"29",x"89",x"3A",x"29",x"2E",x"86",x"CC",x"24",x"6B",x"97",x"B2",x"59",x"55",x"95",x"A8",x"5D",x"CA",x"E9",x"93",x"45",x"3C",x"4E",x"AB",x"9A",x"53",x"75",x"95",x"34",x"25",x"CF",x"C1",x"D4",x"D5",x"9C",x"96",x"3C",x"26",x"75",x"37",x"4B",x"5A",x"D2",x"98",x"35",x"DC",x"B4",x"49",x"8B",x"63",x"F6",x"74",x"D7",x"26",x"2D",x"CA",x"31",x"52",x"43",x"9B",x"B4",x"28",x"7B",x"4D",x"73",x"6F",x"DA",x"92",x"EA",x"CC",x"CD",x"AC",x"6E",x"4B",x"BA",x"0B",x"31",x"D5",x"39",x"23",x"99",x"B6",x"84",x"5D",x"17",x"8F",x"64",x"FA",x"61",x"2C",x"AD",x"D5",x"D2",x"EE",x"9D",x"B2",x"A8",x"EC",x"48",x"5A",x"30",x"F1",x"A4",x"AA",x"23",x"AA",x"51",x"DD",x"2C",x"6B",x"8F",x"B0",x"14",x"B7",x"D0",x"AA",x"32",x"A2",x"DC",x"52",x"D2",x"AB",x"EC",x"88",x"73",x"4D",x"0F",x"AB",x"2A",x"23",x"CE",x"35",x"DD",x"AD",x"EB",x"8C",x"24",x"D5",x"72",x"8B",x"9C",x"32",x"D2",x"14",x"AB",x"9C",x"B3",x"C9",x"C8",x"93",x"AD",x"4A",x"F2",x"26",x"AD",x"4C",x"2E",x"32",x"D8",x"63",x"B7",x"2A",x"79",x"8F",x"10",x"B7",x"D4",x"DA",x"9C",x"DC",x"4C",x"D3",x"36",x"01",x"4A",x"2E",x"77",x"71",x"2E",x"15",x"66",x"5D",x"D7",x"A5",x"45",x"4F",x"A4",x"D8",x"12",x"91",x"55",x"5E",x"31",x"CA",x"4D",x"09",x"D0",x"65",x"D8",x"03",x"FF",
		x"60",x"04",x"98",x"3C",x"0D",x"01",x"C5",x"86",x"B7",x"B8",x"F8",x"0C",x"8B",x"AC",x"33",x"C2",x"62",x"36",x"2C",x"62",x"F6",x"08",x"8A",x"DA",x"F4",x"F0",x"D9",x"23",x"2C",x"66",x"D2",x"C3",x"27",x"8F",x"A8",x"B8",x"09",x"0B",x"9F",x"32",x"E2",x"E6",x"37",x"CD",x"6D",x"F6",x"48",x"5A",x"1A",x"57",x"B3",x"39",x"23",x"ED",x"A5",x"5C",x"D4",x"9B",x"8C",x"B4",x"67",x"53",x"B5",x"8C",x"32",x"D2",x"91",x"9C",x"4D",x"32",x"EA",x"C8",x"9A",x"37",x"33",x"89",x"A8",x"23",x"AB",x"BE",x"5C",x"54",x"2B",x"8F",x"AC",x"C5",x"50",x"51",x"AB",x"32",x"F2",x"E6",x"4D",x"D8",x"A3",x"76",x"AB",x"7A",x"54",x"11",x"CD",x"38",x"AD",x"E9",x"21",x"D8",x"C4",x"EB",x"B4",x"AE",x"EB",x"60",x"17",x"6F",x"D2",x"8A",x"14",x"CD",x"D5",x"BA",x"6E",x"AB",x"92",x"AD",x"0C",x"8E",x"A9",x"AD",x"CA",x"7A",x"32",x"44",x"E7",x"B4",x"BA",x"E8",x"AE",x"12",x"99",x"D3",x"AA",x"6C",x"A7",x"5C",x"74",x"4A",x"AB",x"8B",x"EF",x"34",x"D1",x"3A",x"AD",x"AE",x"C9",x"8A",x"C9",x"9C",x"B6",x"A6",x"64",x"0F",x"E2",x"B4",x"D3",x"9A",x"A2",x"25",x"9C",x"3D",x"6A",x"69",x"8A",x"D2",x"08",x"92",x"B0",x"A5",x"CD",x"46",x"23",x"88",x"EB",x"94",x"26",x"1B",x"37",x"25",x"9E",x"53",x"AA",x"6C",x"3D",x"8D",x"6D",x"4E",x"AB",x"B3",x"8B",x"31",x"C9",x"26",x"AD",x"2E",x"36",x"27",x"C4",x"EB",x"B4",x"BA",x"D8",x"18",x"37",x"AB",x"D3",x"EA",x"EA",x"72",x"DC",x"AD",x"4E",x"6B",x"AA",x"CB",x"76",x"F3",x"25",x"AD",x"AD",x"3E",x"CB",x"DC",x"D7",x"B4",x"B6",x"87",x"74",x"73",x"5B",x"D3",x"BA",x"11",x"D2",x"44",x"6D",x"4E",x"EB",x"A6",x"2B",x"63",x"95",x"C9",x"AD",x"6D",x"AE",x"5C",x"D4",x"2B",x"97",x"A6",x"E9",x"AE",x"54",x"6F",x"9C",x"DA",x"66",x"27",x"43",x"7D",x"89",x"00",x"86",x"69",x"67",x"C0",x"F4",x"ED",x"0C",x"58",x"AE",x"83",x"01",x"5D",x"85",x"A4",x"3E",x"56",x"75",x"A9",x"B1",x"53",x"86",x"14",x"BD",x"71",x"26",x"55",x"99",x"72",x"8C",x"E6",x"E8",x"BA",x"65",x"4E",x"25",x"8A",x"AA",x"13",x"97",x"A5",x"78",x"1F",x"CE",x"6C",x"52",x"96",x"9C",x"BD",x"68",x"AA",x"71",x"59",x"73",x"F3",x"E4",x"9E",x"54",x"69",x"4B",x"4D",x"DD",x"B6",x"92",x"A4",x"AD",x"54",x"77",x"9A",x"98",x"93",x"B6",x"9C",x"34",x"A5",x"2B",x"6A",x"DA",x"8B",x"D1",x"D6",x"F0",x"29",x"69",x"2F",x"51",x"42",x"3A",x"ED",x"84",x"BD",x"3A",x"4D",x"AA",x"A8",x"0A",x"EC",x"28",x"4E",x"5C",x"6A",x"AA",x"A0",x"23",x"69",x"B1",x"E8",x"9D",x"FC",x"00",x"FF",
		x"60",x"04",x"18",x"B5",x"8D",x"01",x"DD",x"B0",x"14",x"BF",x"65",x"36",x"8B",x"A8",x"3D",x"9C",x"5E",x"CA",x"C4",x"75",x"C9",x"30",x"7B",x"1E",x"35",x"F5",x"25",x"C3",x"E8",x"A5",x"CD",x"C5",x"1A",x"0F",x"73",x"84",x"14",x"65",x"5F",x"DC",x"9C",x"AA",x"C8",x"52",x"2B",x"4E",x"F1",x"8A",x"61",x"77",x"8E",x"28",x"C3",x"9F",x"CE",x"45",x"D5",x"6A",x"0F",x"7F",x"F9",x"20",x"B6",x"68",x"3C",x"82",x"5E",x"8A",x"58",x"AD",x"CB",x"08",x"6B",x"34",x"09",x"91",x"36",x"23",x"2E",x"5E",x"22",x"94",x"DB",x"B4",x"AC",x"06",x"B6",x"30",x"49",x"52",x"B2",x"16",x"49",x"D2",x"35",x"6E",x"CB",x"9B",x"15",x"8A",x"50",x"67",x"23",x"2B",x"59",x"DD",x"C8",x"DA",x"8C",x"B4",x"95",x"34",x"13",x"6B",x"33",x"92",x"9E",x"D3",x"54",x"A2",x"CD",x"08",x"7B",x"74",x"15",x"EB",x"36",x"C3",x"1F",x"C9",x"94",x"AC",x"9B",x"34",x"BF",x"07",x"26",x"E9",x"6E",x"12",x"BC",x"9E",x"59",x"4D",x"D5",x"09",x"01",x"84",x"94",x"66",x"40",x"37",x"C4",x"C5",x"6A",x"81",x"D8",x"B3",x"9B",x"36",x"B3",x"58",x"D6",x"CC",x"6E",x"D2",x"8C",x"E2",x"44",x"23",x"26",x"49",x"33",x"8B",x"17",x"B1",x"18",x"27",x"CA",x"CD",x"8E",x"2D",x"7A",x"E4",x"02",x"02",x"16",x"09",x"53",x"46",x"33",x"CA",x"9E",x"95",x"C4",x"18",x"5D",x"07",x"99",x"E7",x"12",x"61",x"36",x"E3",x"6C",x"56",x"75",x"11",x"90",x"A4",x"E9",x"03",x"FF",
		x"60",x"0C",x"38",x"B5",x"53",x"00",x"DD",x"90",x"36",x"BB",x"18",x"63",x"CB",x"58",x"33",x"EC",x"E4",x"2D",x"2C",x"A2",x"D1",x"70",x"92",x"2D",x"37",x"EF",x"D4",x"C3",x"C9",x"B6",x"22",x"A4",x"5A",x"0F",x"37",x"DB",x"8E",x"90",x"6E",x"3C",x"DC",x"62",x"CA",x"83",x"BA",x"4E",x"F3",x"8B",x"4B",x"53",x"DC",x"24",x"04",x"98",x"24",x"84",x"00",x"87",x"BB",x"39",x"A7",x"98",x"8E",x"E0",x"6C",x"EC",x"DC",x"A2",x"3B",x"42",x"B3",x"B5",x"73",x"AB",x"1C",x"0B",x"AE",x"26",x"CE",x"2F",x"A6",x"D4",x"69",x"EB",x"00",x"30",x"60",x"78",x"51",x"06",x"6C",x"6D",x"2C",x"80",x"15",x"55",x"19",x"30",x"B4",x"59",x"1B",x"67",x"D3",x"20",x"B3",x"75",x"6D",x"9C",x"45",x"82",x"DC",x"B6",x"B5",x"71",x"16",x"2B",x"32",x"DD",x"DA",x"C6",x"91",x"AD",x"C8",x"6C",x"2B",x"1B",x"46",x"F6",x"66",x"A1",x"AD",x"6D",x"EA",x"D1",x"0A",x"CC",x"9E",x"B6",x"A9",x"27",x"4D",x"B0",x"5C",x"DB",x"C6",x"11",x"35",x"50",x"E3",x"5D",x"9B",x"46",x"F1",x"24",x"D1",x"65",x"6D",x"9A",x"C5",x"83",x"44",x"97",x"B6",x"79",x"64",x"57",x"32",x"9B",x"D3",x"E6",x"9E",x"44",x"39",x"AC",x"6E",x"9B",x"7B",x"92",x"20",x"B3",x"26",x"6D",x"EE",x"81",x"9D",x"C2",x"EA",x"B4",x"A5",x"07",x"76",x"0A",x"AF",x"5A",x"D6",x"11",x"C5",x"44",x"A4",x"6A",x"5A",x"9B",x"17",x"95",x"B0",x"28",x"6E",x"6B",x"8E",x"CC",x"D3",x"A2",x"3C",x"FF",
		x"60",x"08",x"28",x"2A",x"1D",x"01",x"D5",x"84",x"13",x"A0",x"59",x"F7",x"50",x"86",x"E4",x"69",x"AC",x"4D",x"4A",x"E5",x"7D",x"86",x"B2",x"B4",x"69",x"79",x"D0",x"99",x"C9",x"DC",x"A5",x"45",x"51",x"57",x"26",x"72",x"97",x"E6",x"47",x"59",x"55",x"84",x"9D",x"8B",x"EB",x"D4",x"76",x"0A",x"B7",x"4E",x"76",x"60",x"3B",x"AE",x"D2",x"26",x"19",x"09",x"CD",x"8A",x"6A",x"DB",x"E0",x"14",x"92",x"E9",x"24",x"6D",x"95",x"57",x"78",x"44",x"86",x"5A",x"6E",x"F9",x"52",x"CE",x"2A",x"DE",x"75",x"E4",x"8D",x"0B",x"47",x"56",x"AB",x"51",x"74",x"AB",x"64",x"9E",x"9D",x"46",x"5E",x"A3",x"B0",x"69",x"75",x"19",x"59",x"09",x"22",x"66",x"D1",x"A5",x"65",x"D9",x"1B",x"87",x"E4",x"D6",x"92",x"67",x"AF",x"1E",x"EC",x"5D",x"42",x"16",x"9D",x"7A",x"B2",x"77",x"51",x"49",x"74",x"D2",x"AE",x"D6",x"55",x"C5",x"C9",x"89",x"A5",x"67",x"2D",x"95",x"25",x"6F",x"12",x"92",x"9B",x"59",x"9E",x"BC",x"5A",x"B0",x"77",x"21",x"59",x"74",x"1A",x"C1",x"DE",x"85",x"A4",x"C1",x"69",x"86",x"58",x"97",x"07",x"FF",
		x"60",x"61",x"19",x"01",x"4A",x"D9",x"F3",x"96",x"A9",x"6A",x"2E",x"45",x"EB",x"DA",x"BA",x"62",x"AC",x"5C",x"BC",x"5B",x"6B",x"92",x"B1",x"0A",x"93",x"AD",x"AD",x"A9",x"4A",x"B3",x"8C",x"B5",x"B9",x"3A",x"59",x"2D",x"13",x"4D",x"03",x"02",x"C8",x"A3",x"51",x"01",x"D5",x"96",x"29",x"A0",x"CB",x"31",x"05",x"74",x"11",x"82",x"01",x"D7",x"39",x"5B",x"5E",x"24",x"6D",x"4B",x"E7",x"DC",x"24",x"73",x"D4",x"69",x"6D",x"52",x"B9",x"C2",x"D1",x"B8",x"B5",x"55",x"E9",x"A9",x"DB",x"9A",x"D6",x"36",x"63",x"6B",x"6E",x"AB",x"5B",x"DB",x"6C",x"B4",x"84",x"2D",x"6B",x"4D",x"8D",x"E1",x"E2",x"39",x"37",x"34",x"23",x"A4",x"30",x"C7",x"52",x"02",x"44",x"C6",x"A9",x"DA",x"24",x"B3",x"9D",x"DC",x"AE",x"6B",x"AB",x"D2",x"33",x"B7",x"D6",x"A1",x"6D",x"DA",x"36",x"D4",x"DB",x"10",x"20",x"10",x"E9",x"54",x"76",x"17",x"2E",x"A2",x"49",x"5A",x"D9",x"8A",x"13",x"6B",x"B4",x"6B",x"79",x"8D",x"CA",x"A6",x"96",x"AD",x"65",x"D9",x"04",x"BB",x"68",x"BA",x"92",x"24",x"59",x"E2",x"8E",x"ED",x"52",x"E2",x"6D",x"B8",x"8B",x"37",x"49",x"69",x"CC",x"26",x"EA",x"16",x"B7",x"65",x"59",x"A4",x"49",x"50",x"BA",x"96",x"55",x"6C",x"AE",x"CD",x"69",x"5A",x"5C",x"94",x"9B",x"2B",x"D5",x"69",x"61",x"56",x"A1",x"E6",x"B2",x"B8",x"F9",x"49",x"BB",x"78",x"E8",x"92",x"E6",x"25",x"E3",x"12",x"A1",x"4B",x"9B",x"97",x"8C",x"4B",x"B8",x"2C",x"6D",x"5E",x"B2",x"A6",x"A1",x"BA",x"AE",x"F9",x"D1",x"8B",x"07",x"5B",x"B7",x"16",x"44",x"A7",x"11",x"AA",x"ED",x"5A",x"18",x"9D",x"46",x"1A",x"B7",x"6B",x"49",x"08",x"EE",x"26",x"DC",x"B6",x"A5",x"D1",x"67",x"AA",x"62",x"B2",x"96",x"05",x"E3",x"19",x"CA",x"C9",x"5A",x"1E",x"AC",x"47",x"1A",x"A5",x"6D",x"79",x"70",x"16",x"A6",x"9A",x"B6",x"E5",x"D1",x"59",x"98",x"69",x"D3",x"52",x"64",x"ED",x"26",x"66",x"4D",x"53",x"DD",x"B9",x"8B",x"07",x"A7",x"61",x"40",x"63",x"19",x"26",x"1B",x"CC",x"AD",x"82",x"6D",x"9B",x"6C",x"13",x"73",x"4D",x"93",x"A3",x"B2",x"C9",x"CC",x"35",x"D9",x"35",x"CB",x"33",x"4B",x"75",x"53",x"B7",x"08",x"A8",x"54",x"E4",x"01",x"FF",
		x"60",x"0C",x"A8",x"49",x"42",x"00",x"AD",x"46",x"0A",x"A0",x"B4",x"F4",x"64",x"A5",x"2A",x"A9",x"A5",x"93",x"87",x"59",x"B2",x"9B",x"A5",x"AD",x"1E",x"56",x"8D",x"21",x"9E",x"B1",x"64",x"D8",x"2D",x"A9",x"AA",x"D7",x"94",x"E6",x"B5",x"48",x"C2",x"5D",x"55",x"52",x"B4",x"D6",x"84",x"28",x"A9",x"56",x"C0",x"AC",x"AE",x"0A",x"E8",x"49",x"A2",x"A5",x"B5",x"89",x"68",x"F8",x"92",x"96",x"E5",x"4C",x"A6",x"19",x"CD",x"5A",x"95",x"07",x"69",x"84",x"B6",x"6B",x"5D",x"1E",x"2A",x"92",x"9E",x"BC",x"0D",x"B9",x"A9",x"48",x"7A",x"F2",x"36",x"E5",x"C5",x"2E",x"EE",x"F1",x"C2",x"92",x"0F",x"B9",x"BB",x"2C",x"61",x"7B",x"DE",x"18",x"61",x"BE",x"13",x"1D",x"B9",x"A3",x"8D",x"45",x"4A",x"00",x"10",x"83",x"91",x"5B",x"A1",x"62",x"45",x"D5",x"52",x"6F",x"BA",x"4A",x"65",x"97",x"1B",x"B5",x"15",x"46",x"B3",x"5B",x"E2",x"ED",x"97",x"B2",x"2C",x"1E",x"41",x"B4",x"57",x"62",x"B6",x"64",x"78",x"29",x"8D",x"AB",x"E5",x"94",x"E1",x"E6",x"E0",x"2E",x"5E",x"51",x"82",x"13",x"0C",x"87",x"64",x"DA",x"4E",x"5E",x"32",x"12",x"5C",x"E5",x"AA",x"84",x"D1",x"85",x"7A",x"A7",x"98",x"11",x"E4",x"D0",x"6E",x"15",x"66",x"5A",x"90",x"5D",x"99",x"94",x"55",x"19",x"7E",x"CE",x"6E",x"92",x"51",x"B6",x"F9",x"C5",x"6B",x"92",x"65",x"1C",x"E5",x"65",x"8F",x"C1",x"99",x"69",x"4A",x"50",x"26",x"07",x"B9",x"B7",x"6E",x"41",x"CE",x"94",x"66",x"B2",x"28",x"05",x"31",x"53",x"99",x"C6",x"AC",x"12",x"E6",x"84",x"A5",x"9E",x"B3",x"8D",x"5F",x"22",x"A5",x"45",x"35",x"56",x"41",x"A9",x"EC",x"62",x"D6",x"5A",x"04",x"29",x"73",x"04",x"5B",x"2B",x"11",x"A4",x"4C",x"9E",x"E2",x"AD",x"00",x"01",x"4E",x"8B",x"BA",x"AC",x"88",x"A8",x"4A",x"8C",x"13",x"12",x"B7",x"CB",x"C4",x"A3",x"4A",x"4A",x"7C",x"99",x"14",x"B3",x"26",x"2D",x"4B",x"6E",x"D2",x"4C",x"1B",x"B7",x"A2",x"86",x"74",x"53",x"6D",x"DC",x"DA",x"5E",x"52",x"44",x"A2",x"76",x"9A",x"46",x"0C",x"12",x"AB",x"D1",x"00",x"04",x"28",x"3A",x"8D",x"00",x"8B",x"A6",x"21",x"E0",x"C9",x"36",x"04",x"1C",x"59",x"8A",x"80",x"23",x"DA",x"11",x"B0",x"79",x"FB",x"03",x"FF",
		x"60",x"2B",x"E8",x"32",x"CC",x"CD",x"6C",x"EF",x"60",x"07",x"3B",x"D8",x"C1",x"0E",x"76",x"B0",x"83",x"1D",x"EC",x"60",x"07",x"3B",x"D8",x"C1",x"0E",x"76",x"B0",x"83",x"1D",x"EC",x"60",x"07",x"3B",x"D8",x"C1",x"0E",x"76",x"B0",x"83",x"1D",x"EC",x"60",x"07",x"3B",x"D8",x"C1",x"0E",x"76",x"B0",x"83",x"1D",x"EC",x"60",x"07",x"3B",x"D8",x"C1",x"0E",x"76",x"B0",x"83",x"07",x"FF",
		x"60",x"AD",x"4E",x"56",x"DD",x"32",x"AC",x"B4",x"2A",x"65",x"35",x"AD",x"A8",x"DA",x"B2",x"E4",x"A3",x"55",x"A5",x"4D",x"4B",x"93",x"F2",x"35",x"A5",x"34",x"2D",x"08",x"36",x"57",x"D4",x"1C",x"37",x"3F",x"38",x"6B",x"11",x"57",x"93",x"BC",x"E0",x"D5",x"D4",x"CA",x"B2",x"02",x"6A",x"08",x"45",x"C0",x"70",x"69",x"04",x"98",x"AD",x"9C",x"01",x"A3",x"B5",x"0B",x"A0",x"F7",x"EA",x"96",x"E5",x"28",x"A2",x"EE",x"AD",x"47",x"55",x"2C",x"85",x"9A",x"F6",x"1E",x"6D",x"B1",x"A2",x"22",x"91",x"96",x"01",x"B3",x"A6",x"22",x"A0",x"39",x"66",x"04",x"D4",x"2A",x"52",x"FA",x"E4",x"9D",x"D2",x"7B",x"CA",x"E8",x"92",x"77",x"75",x"89",x"39",x"A6",x"4D",x"DC",x"55",x"D3",x"6B",x"03",x"30",x"20",x"58",x"E6",x"56",x"55",x"5D",x"1E",x"6A",x"51",x"5A",x"9D",x"6D",x"46",x"92",x"97",x"69",x"AD",x"6F",x"ED",x"62",x"39",x"7B",x"34",x"DE",x"77",x"3A",x"D9",x"9A",x"51",x"FA",x"30",x"A1",x"EC",x"AD",x"47",x"EA",x"62",x"86",x"52",x"AC",x"4E",x"71",x"A8",x"A6",x"2C",x"51",x"9B",x"01",x"75",x"57",x"29",x"A0",x"F5",x"4E",x"03",x"B4",x"31",x"25",x"80",x"76",x"2A",x"47",x"97",x"3D",x"B9",x"8D",x"C7",x"1A",x"6D",x"A9",x"22",x"9A",x"D5",x"64",x"0C",x"2D",x"A6",x"8B",x"C4",x"92",x"D1",x"B5",x"E0",x"29",x"14",x"89",x"47",x"55",x"0C",x"8B",x"DA",x"A8",x"6E",x"49",x"B6",x"EC",x"54",x"E1",x"B2",x"05",x"C9",x"B1",x"6A",x"94",x"CA",x"E6",x"67",x"2F",x"86",x"9D",x"B1",x"4B",x"58",x"B2",x"09",x"46",x"C7",x"76",x"59",x"C9",x"2E",x"48",x"1D",x"CB",x"14",x"59",x"8A",x"9B",x"8C",x"22",x"15",x"65",x"65",x"2A",x"1E",x"B1",x"85",x"1F",x"95",x"A9",x"59",x"3B",x"64",x"41",x"36",x"A6",x"E2",x"1D",x"8B",x"C4",x"C5",x"AA",x"92",x"77",x"A8",x"07",x"FF",
		x"60",x"2C",x"F0",x"54",x"A3",x"DA",x"12",x"AB",x"94",x"A9",x"9A",x"4E",x"8F",x"A4",x"32",x"CD",x"BD",x"6B",x"C2",x"96",x"CA",x"3D",x"91",x"A9",x"CE",x"C8",x"26",x"D7",x"DC",x"BB",x"C6",x"ED",x"A4",x"2C",x"31",x"8A",x"BA",x"28",x"DD",x"B2",x"A2",x"59",x"FD",x"B2",x"C8",x"C8",x"8A",x"17",x"D7",x"C9",x"22",x"23",x"2D",x"CE",x"83",x"23",x"86",x"8C",x"28",x"C5",x"08",x"AE",x"2C",x"3A",x"FC",x"14",x"32",x"B1",x"32",x"EC",x"70",x"62",x"C8",x"A4",x"CE",x"B0",x"CD",x"0C",x"25",x"8D",x"D6",x"C2",x"36",x"23",x"E4",x"72",x"1C",x"B3",x"DA",x"AC",x"E8",x"3B",x"A1",x"BC",x"58",x"F1",x"82",x"2B",x"C7",x"12",x"3B",x"29",x"B0",x"36",x"82",x"3D",x"A2",x"86",x"48",x"DA",x"08",x"AD",x"88",x"12",x"62",x"61",x"2A",x"AC",x"BC",x"76",x"48",x"98",x"AD",x"8A",x"88",x"3A",x"26",x"65",x"36",x"CA",x"AB",x"AA",x"9A",x"0C",x"C7",x"88",x"AC",x"8E",x"6D",x"0A",x"1C",x"CA",x"B3",x"2B",x"92",x"A9",x"B8",x"75",x"8F",x"EC",x"48",x"A6",x"E2",x"CE",x"C2",x"6B",x"62",x"AB",x"CA",x"5B",x"31",x"AD",x"8E",x"43",x"6A",x"23",x"3C",x"3C",x"2A",x"F6",x"03",x"FF",
		x"60",x"CD",x"2B",x"29",x"3D",x"D6",x"2A",x"37",x"2F",x"A7",x"F4",x"58",x"8D",x"32",x"DC",x"EC",x"27",x"6D",x"24",x"4A",x"73",x"52",x"A9",x"8C",x"D5",x"C0",x"4D",x"4F",x"23",x"22",x"5A",x"AB",x"0C",x"25",x"8D",x"8A",x"E8",x"2C",x"D3",x"E4",x"78",x"33",x"AD",x"2A",x"72",x"93",x"E3",x"8D",x"94",x"6E",x"CB",x"4D",x"8D",x"3B",x"8B",x"2A",x"23",x"15",x"3D",x"EC",x"2C",x"AA",x"AC",x"D5",x"9C",x"30",x"B3",x"20",x"72",x"56",x"F1",x"7D",x"AF",x"82",x"8C",x"D9",x"29",x"74",x"37",x"0C",x"AB",x"E3",x"A4",x"58",x"F7",x"0E",x"B4",x"4E",x"92",x"52",x"99",x"BB",x"99",x"33",x"A9",x"CB",x"78",x"9F",x"42",x"CD",x"24",x"AA",x"54",x"AE",x"97",x"D8",x"93",x"D0",x"FA",x"01",x"FF",
		x"60",x"C3",x"6D",x"B6",x"5B",x"B3",x"EA",x"0E",x"37",x"E7",x"72",x"DB",x"8A",x"32",x"AC",x"94",x"A7",x"A4",x"23",x"EA",x"50",x"73",x"98",x"D6",x"AC",x"44",x"43",x"49",x"B9",x"8B",x"3D",x"1A",x"0F",x"35",x"D6",x"74",x"4E",x"AF",x"3D",x"8C",x"30",x"83",x"A9",x"BC",x"49",x"71",x"43",x"70",x"17",x"CB",x"73",x"25",x"2C",x"C6",x"C3",x"04",x"1F",x"9B",x"28",x"1B",x"49",x"37",x"59",x"82",x"00",x"5D",x"45",x"40",x"00",x"C3",x"48",x"30",x"E0",x"78",x"53",x"01",x"6C",x"EF",x"A1",x"80",x"9D",x"22",x"15",x"B0",x"82",x"BB",x"02",x"66",x"CA",x"10",x"C0",x"48",x"19",x"04",x"E8",x"5E",x"15",x"01",x"55",x"90",x"3E",x"FF",
		x"60",x"45",x"4C",x"B6",x"1A",x"DD",x"AF",x"35",x"CE",x"97",x"0C",x"9A",x"8A",x"D2",x"58",x"1F",x"32",x"29",x"32",x"4C",x"11",x"4C",x"C8",x"C4",x"C8",x"50",x"49",x"D6",x"25",x"43",x"A2",x"22",x"25",x"55",x"D7",x"08",x"A9",x"AE",x"98",x"0C",x"97",x"DC",x"B9",x"62",x"B6",x"73",x"5D",x"8C",x"E0",x"88",x"99",x"2E",x"08",x"26",x"8B",x"52",x"67",x"AA",x"38",x"04",x"37",x"72",x"9F",x"45",x"93",x"07",x"FF",
		x"60",x"41",x"28",x"3C",x"D6",x"4C",x"EB",x"16",x"DE",x"DB",x"5E",x"35",x"9F",x"5A",x"F8",x"10",x"A6",x"D1",x"63",x"6C",x"E1",x"42",x"E9",x"82",x"AC",x"A8",x"89",x"F3",x"B9",x"13",x"3C",x"83",x"25",x"DE",x"E7",x"0E",x"88",x"AC",x"5C",x"04",x"97",x"3B",x"20",x"32",x"71",x"92",x"5C",x"E8",x"02",x"0B",x"37",x"41",x"15",x"A5",x"13",x"3C",x"1C",x"3B",x"4B",x"84",x"1E",x"C8",x"8C",x"69",x"5C",x"91",x"DB",x"49",x"22",x"89",x"0A",x"85",x"9D",x"16",x"F6",x"BA",x"22",x"55",x"A2",x"CB",x"4D",x"AD",x"D2",x"EC",x"01",x"FF",
		x"60",x"4C",x"D4",x"B5",x"43",x"C8",x"9D",x"28",x"81",x"E7",x"0E",x"13",x"B3",x"63",x"78",x"D6",x"52",x"CD",x"32",x"49",x"E0",x"78",x"0D",x"35",x"F7",x"B8",x"81",x"E3",x"39",x"4D",x"22",x"ED",x"05",x"8E",x"97",x"54",x"77",x"8F",x"1B",x"58",x"DE",x"5C",x"3D",x"3C",x"69",x"60",x"59",x"0B",x"F1",x"88",x"A4",x"81",x"E3",x"B9",x"C4",x"C2",x"EB",x"05",x"9E",x"55",x"57",x"73",x"4F",x"EA",x"04",x"D6",x"5C",x"CC",x"3D",x"A9",x"51",x"79",x"4B",x"11",x"B5",x"24",x"4A",x"67",x"B9",x"55",x"45",x"93",x"30",x"9B",x"85",x"09",x"57",x"B1",x"C3",x"7C",x"A9",x"3A",x"33",x"4D",x"0E",x"0A",x"94",x"88",x"EC",x"76",x"D9",x"0F",x"FF",
		x"60",x"C3",x"2D",x"B1",x"D2",x"36",x"9A",x"0C",x"2B",x"CD",x"88",x"5C",x"B3",x"32",x"F4",x"34",x"3D",x"7D",x"35",x"CA",x"50",x"D3",x"F2",x"88",x"D5",x"C4",x"43",x"8E",x"37",x"3D",x"C6",x"42",x"0F",x"31",x"8D",x"09",x"6D",x"2B",x"D2",x"C4",x"78",x"D3",x"35",x"33",x"4C",x"11",x"E2",x"73",x"D3",x"4E",x"2B",x"41",x"0C",x"DF",x"43",x"AA",x"CD",x"24",x"29",x"EC",x"4C",x"CA",x"2C",x"55",x"D4",x"70",x"23",x"B0",x"2A",x"72",x"32",x"FD",x"09",x"A7",x"4A",x"CB",x"C1",x"F5",x"BD",x"12",x"A2",x"62",x"B9",x"C0",x"8D",x"76",x"F0",x"6A",x"62",x"22",x"73",x"53",x"38",x"A6",x"A9",x"4A",x"D4",x"2A",x"43",x"EF",x"26",x"22",x"D5",x"79",x"0A",x"B9",x"92",x"D0",x"FC",x"01",x"FF",
		x"60",x"CA",x"1D",x"86",x"18",x"27",x"AA",x"2A",x"37",x"11",x"89",x"5C",x"B1",x"E2",x"B4",x"28",x"D9",x"7B",x"38",x"4A",x"93",x"82",x"D1",x"AE",x"55",x"BB",x"43",x"AE",x"49",x"DD",x"26",x"CC",x"0D",x"29",x"67",x"2D",x"EF",x"34",x"3F",x"E4",x"5C",x"BC",x"ED",x"DC",x"CA",x"90",x"F2",x"8C",x"B4",x"0E",x"AB",x"43",x"89",x"BD",x"C2",x"DA",x"A3",x"16",x"39",x"CE",x"4E",x"EE",x"A8",x"5A",x"E4",x"B0",x"BA",x"B0",x"B3",x"6A",x"D1",x"C2",x"EC",x"C6",x"88",x"31",x"C9",x"F2",x"6B",x"1A",x"C2",x"AA",x"24",x"C7",x"8F",x"69",x"C8",x"A8",x"95",x"3C",x"DF",x"66",x"C0",x"B2",x"76",x"F0",x"6D",x"9D",x"01",x"8D",x"5A",x"2E",x"D4",x"A5",x"07",x"BC",x"6A",x"9B",x"48",x"9C",x"76",x"F4",x"B4",x"A3",x"62",x"99",x"A6",x"51",x"22",x"89",x"48",x"AC",x"CA",x"75",x"56",x"3B",x"34",x"7F",x"FF",
		x"60",x"CD",x"8F",x"A3",x"42",x"26",x"A3",x"0E",x"2F",x"D5",x"4E",x"9E",x"0C",x"33",x"BC",x"D4",x"3A",x"64",x"22",x"EC",x"70",x"53",x"E8",x"E6",x"8A",x"B0",x"C3",x"49",x"61",x"9A",x"2B",x"C2",x"0E",x"3B",x"85",x"69",x"CE",x"0C",x"3B",x"9C",x"14",x"A6",x"39",x"B3",x"EC",x"70",x"B3",x"9F",x"A6",x"8C",x"30",x"C3",x"CB",x"6E",x"9A",x"2A",x"A2",x"0C",x"2F",x"96",x"09",x"29",x"0F",x"3D",x"FC",x"C6",x"63",x"34",x"D5",x"F4",x"08",x"8A",x"EE",x"D6",x"90",x"C2",x"2D",x"2C",x"BA",x"4A",x"4D",x"4B",x"B7",x"A8",x"98",x"6A",x"33",x"2D",x"54",x"E2",x"AA",x"B2",x"D4",x"A5",x"70",x"49",x"8B",x"CB",x"56",x"B3",x"D2",x"25",x"2F",x"A6",x"5B",x"CA",x"82",x"AA",x"A2",x"2A",x"5F",x"13",x"29",x"FC",x"00",x"FF",
		x"60",x"CD",x"48",x"AE",x"56",x"4C",x"C7",x"36",x"3D",x"B9",x"5A",x"31",x"9D",x"DB",x"CC",x"10",x"7B",x"38",x"6C",x"6E",x"33",x"42",x"EE",x"C2",x"B0",x"2A",x"4D",x"0D",x"B9",x"0B",x"D2",x"CA",x"34",x"25",x"9A",x"1E",x"48",x"9B",x"DA",x"A4",x"68",x"6B",x"51",x"7D",x"4C",x"91",x"A3",x"ED",x"45",x"F5",x"31",x"45",x"89",x"A6",x"97",x"44",x"87",x"14",x"25",x"84",x"19",x"30",x"AF",x"5C",x"B4",x"E0",x"7A",x"51",x"BD",x"72",x"D2",x"7D",x"9E",x"86",x"F0",x"B2",x"49",x"B3",x"79",x"0A",x"C2",x"CB",x"26",x"C3",x"BB",x"19",x"30",x"2F",x"92",x"4C",x"EF",x"67",x"C0",x"7C",x"74",x"B2",x"BD",x"A9",x"45",x"B5",x"C9",x"C1",x"75",x"7E",x"06",x"CC",x"6B",x"39",x"3F",x"A8",x"3C",x"12",x"9D",x"65",x"42",x"AF",x"F2",x"88",x"75",x"B6",x"89",x"BC",x"AE",x"23",x"D6",x"DA",x"2E",x"F1",x"3A",x"97",x"58",x"E3",x"A8",x"D4",x"B8",x"1E",x"64",x"4B",x"FA",x"00",x"FF",
		x"60",x"86",x"35",x"B3",x"9C",x"39",x"92",x"26",x"56",x"AF",x"72",x"D6",x"88",x"94",x"18",x"B3",x"2A",x"C9",x"B4",x"72",x"A2",x"4D",x"EF",x"22",x"E5",x"D8",x"89",x"31",x"6D",x"8A",x"94",x"9C",x"24",x"C6",x"FA",x"19",x"30",x"56",x"92",x"18",x"ED",x"A7",x"C8",x"2D",x"4E",x"62",x"9D",x"E9",x"46",x"93",x"BA",x"89",x"93",x"B6",x"0B",x"53",x"93",x"06",x"5E",x"E6",x"4A",x"08",x"AB",x"9B",x"44",x"ED",x"A6",x"21",x"35",x"76",x"92",x"65",x"AE",x"64",x"71",x"27",x"49",x"95",x"B1",x"8B",x"24",x"12",x"27",x"53",x"86",x"6E",x"D2",x"48",x"94",x"6C",x"6D",x"73",x"59",x"6D",x"65",x"72",x"44",x"C9",x"20",x"8F",x"DA",x"C1",x"13",x"AE",x"DA",x"DC",x"E4",x"06",x"8F",x"BB",x"CC",x"48",x"97",x"1D",x"22",x"EB",x"DC",x"3D",x"D5",x"B2",x"49",x"B8",x"AF",x"74",x"31",x"27",x"0F",x"FF",
		x"60",x"46",x"4E",x"21",x"0B",x"23",x"C7",x"26",x"25",x"C7",x"2A",x"0E",x"1F",x"DB",x"B4",x"EC",x"B3",x"D9",x"A3",x"6C",x"D3",x"52",x"CE",x"E2",x"4A",x"AB",x"4D",x"8D",x"2D",x"42",x"3A",x"AD",x"35",x"35",x"F6",x"70",x"E9",x"B2",x"D6",x"D4",x"D0",x"C3",x"65",x"4A",x"6A",x"53",x"C3",x"74",x"D7",x"29",x"69",x"45",x"0B",x"3D",x"92",x"A7",x"C4",x"16",x"2D",x"94",x"4C",x"EA",x"36",x"DA",x"B4",x"50",x"32",x"39",x"CB",x"6C",x"D1",x"42",x"AD",x"10",x"2F",x"A3",x"45",x"F7",x"B5",x"52",x"BC",x"8D",x"34",x"2B",x"94",x"0C",x"C9",x"0E",x"D3",x"EC",x"90",x"33",x"B9",x"2A",x"CC",x"70",x"62",x"CC",x"E4",x"E8",x"28",x"C3",x"8D",x"31",x"8B",x"A3",x"C2",x"0C",x"37",x"FA",x"2C",x"B1",x"2A",x"DD",x"BC",x"90",x"A2",x"A8",x"3A",x"74",x"F1",x"43",x"B3",x"A0",x"E9",x"30",x"25",x"0C",x"D5",x"82",x"A7",x"43",x"A7",x"28",x"E4",x"08",x"AD",x"2C",x"12",x"92",x"90",x"D5",x"6D",x"C2",x"48",x"48",x"73",x"31",x"A3",x"88",x"B0",x"2C",x"CD",x"DE",x"8C",x"34",x"2A",x"3D",x"FF",
		x"60",x"C9",x"48",x"BE",x"8A",x"3D",x"C7",x"24",x"2D",x"E6",x"4E",x"8A",x"1A",x"92",x"94",x"38",x"43",x"65",x"CA",x"48",x"91",x"43",x"2F",x"93",x"C9",x"20",x"4D",x"8E",x"BE",x"8B",x"3D",x"07",x"37",x"39",x"E6",x"4A",x"CA",x"2E",x"DC",x"E4",x"98",x"2B",x"39",x"BA",x"48",x"93",x"63",x"6E",x"E7",x"AA",x"22",x"4D",x"8E",x"A5",x"9C",x"B3",x"0B",x"37",x"39",x"96",x"36",x"EE",x"2E",x"52",x"E4",x"58",x"CB",x"78",x"AA",x"48",x"51",x"62",x"2D",x"A7",x"EE",x"C2",x"45",x"8D",x"B9",x"83",x"B2",x"87",x"14",x"35",x"A6",x"4A",x"8A",x"1E",x"53",x"B4",x"98",x"3B",x"A8",x"6A",x"6C",x"D1",x"63",x"EE",x"A0",x"AA",x"71",x"C5",x"88",x"B1",x"93",x"A2",x"86",x"17",x"23",x"C6",x"2A",x"8A",x"1A",x"56",x"CC",x"50",x"CA",x"B9",x"7A",x"6C",x"B1",x"62",x"A9",x"A0",x"EA",x"B1",x"C5",x"8E",x"B9",x"12",x"73",x"C6",x"14",x"27",x"A6",x"2A",x"8C",x"19",x"53",x"DC",x"18",x"AB",x"30",x"7A",x"4C",x"71",x"A3",x"AF",x"22",x"CB",x"33",x"C5",x"8B",x"3E",x"9B",x"BC",x"A6",x"14",x"2F",x"9A",x"1C",x"D1",x"98",x"5A",x"FC",x"68",x"62",x"CC",x"6C",x"4C",x"F1",x"43",x"C8",x"12",x"8F",x"31",x"C5",x"0F",x"A1",x"52",x"32",x"C6",x"94",x"20",x"86",x"4A",x"F6",x"38",x"53",x"82",x"E4",x"AB",x"C8",x"FC",x"72",x"0A",x"52",x"AC",x"22",x"F3",x"D3",x"29",x"8C",x"B1",x"8A",x"CC",x"2F",x"A7",x"30",x"86",x"2A",x"32",x"BF",x"92",x"C2",x"E8",x"AB",x"C9",x"FC",x"4A",x"8A",x"92",x"CB",x"66",x"B5",x"2B",x"29",x"4A",x"3E",x"87",x"C5",x"AE",x"A4",x"28",x"D9",x"18",x"11",x"BD",x"9D",x"A2",x"64",x"B3",x"55",x"F5",x"76",x"8A",x"93",x"CB",x"16",x"D5",x"DB",x"29",x"4E",x"26",x"5B",x"8C",x"1E",x"A7",x"38",x"E9",x"6C",x"71",x"5A",x"9C",x"92",x"AC",x"B4",x"4D",x"79",x"72",x"4A",x"B2",x"F0",x"16",x"E3",x"D9",x"21",x"49",x"3A",x"13",x"45",x"66",x"BB",x"34",x"99",x"28",x"12",x"2E",x"6D",x"B2",x"62",x"A2",x"48",x"24",x"12",x"01",x"84",x"72",x"47",x"80",x"92",x"11",x"0F",x"FF",
		x"60",x"0A",x"98",x"B1",x"5D",x"00",x"59",x"90",x"B6",x"AA",x"E7",x"0D",x"62",x"6A",x"3F",x"AA",x"11",x"DA",x"49",x"39",x"FD",x"28",x"87",x"08",x"E3",x"94",x"76",x"A3",x"9A",x"44",x"2A",x"8B",x"D3",x"8C",x"7A",x"22",x"E9",x"4E",x"F2",x"DC",x"EA",x"05",x"65",x"C6",x"48",x"49",x"6B",x"07",x"71",x"D5",x"A9",x"90",x"04",x"C8",x"5A",x"85",x"00",x"49",x"A4",x"12",x"20",x"F0",x"29",x"02",x"04",x"3E",x"2E",x"00",x"6F",x"C4",x"46",x"39",x"5C",x"29",x"48",x"6C",x"19",x"C5",x"B2",x"AE",x"A8",x"B1",x"75",x"64",x"CB",x"77",x"20",x"E8",x"96",x"16",x"8F",x"D8",x"86",x"64",x"5D",x"5A",x"D0",x"4B",x"09",x"8A",x"75",x"49",x"7E",x"EB",x"89",x"64",x"BA",x"96",x"00",x"BD",x"8C",x"33",x"20",x"2B",x"65",x"06",x"14",x"A1",x"4C",x"80",x"2C",x"85",x"10",x"90",x"0D",x"31",x"30",x"A0",x"05",x"D3",x"92",x"97",x"8C",x"EE",x"E6",x"6D",x"5A",x"55",x"2A",x"59",x"A9",x"24",x"6D",x"75",x"71",x"25",x"DA",x"A4",x"B6",x"D5",x"25",x"A5",x"68",x"B2",x"BA",x"D1",x"D4",x"1E",x"22",x"CE",x"5E",x"47",x"3B",x"62",x"39",x"8A",x"B5",x"F3",x"2D",x"30",x"A0",x"1C",x"56",x"06",x"94",x"C1",x"D2",x"B2",x"DA",x"BC",x"82",x"2D",x"F1",x"C8",x"8A",x"EA",x"0C",x"E7",x"A5",x"23",x"AB",x"BC",x"23",x"8A",x"BB",x"B4",x"3C",x"AB",x"76",x"6F",x"D8",x"E2",x"CA",x"62",x"5C",x"A2",x"48",x"4E",x"49",x"93",x"4F",x"D1",x"A6",x"2C",x"25",x"49",x"29",x"D8",x"8A",x"BA",x"94",x"38",x"55",x"27",x"2F",x"EA",x"52",x"E2",x"5C",x"1D",x"BD",x"35",x"4D",x"89",x"4B",x"73",x"71",x"93",x"34",x"02",x"D8",x"4A",x"4D",x"00",x"0D",x"97",x"0B",x"60",x"89",x"4A",x"02",x"04",x"53",x"84",x"80",x"90",x"D0",x"4B",x"70",x"BC",x"A7",x"88",x"24",x"6D",x"41",x"36",x"6E",x"99",x"B2",x"76",x"44",x"95",x"46",x"47",x"51",x"E6",x"16",x"26",x"D2",x"6B",x"2A",x"59",x"4B",x"90",x"F0",x"AC",x"B1",x"B4",x"29",x"41",x"C2",x"B3",x"81",x"D2",x"A6",x"04",x"89",x"E7",x"24",x"59",x"98",x"E6",x"15",x"D2",x"19",x"6A",x"E1",x"9A",x"57",x"C8",x"A4",x"99",x"35",x"69",x"FE",x"C0",x"15",x"6A",x"DE",x"24",x"F9",x"49",x"B9",x"B9",x"45",x"D5",x"E4",x"67",x"19",x"E6",x"9E",x"55",x"5A",x"54",x"74",x"9B",x"5A",x"35",x"69",x"61",x"D1",x"1D",x"66",x"31",x"79",x"C4",x"45",x"77",x"B8",x"C7",x"EC",x"91",x"16",x"3D",x"11",x"1E",x"6B",x"46",x"58",x"5D",x"85",x"BB",x"2F",x"1D",x"41",x"F5",x"69",x"9E",x"31",x"67",x"F8",x"2D",x"85",x"68",x"E4",x"D2",x"E2",x"B7",x"12",x"CC",x"D6",x"4B",x"55",x"D2",x"52",x"89",x"48",x"C6",x"6A",x"6D",x"0D",x"65",x"2A",x"D1",x"B4",x"B5",x"39",x"87",x"AA",x"47",x"D3",x"D6",x"57",x"17",x"E2",x"69",x"51",x"CB",x"D8",x"92",x"B1",x"66",x"45",x"0D",x"4B",x"71",x"EA",x"CA",x"2E",x"37",x"EC",x"D5",x"5B",x"08",x"9B",x"94",x"B0",x"37",x"DB",x"AA",x"1C",x"49",x"1E",x"FF",
		x"60",x"08",x"58",x"48",x"9D",x"01",x"1D",x"88",x"09",x"E0",x"08",x"37",x"01",x"1C",x"95",x"3E",x"92",x"A5",x"8D",x"2B",x"39",x"F3",x"08",x"A2",x"4B",x"77",x"AB",x"3A",x"C3",x"CF",x"62",x"C3",x"C3",x"E7",x"0E",x"27",x"B3",x"4D",x"71",x"9F",x"3D",x"AC",x"24",x"DA",x"4D",x"23",x"76",x"33",x"93",x"2A",x"37",x"0A",x"D1",x"C9",x"89",x"B2",x"4D",x"D9",x"2D",x"A5",x"30",x"D9",x"72",x"35",x"8F",x"3D",x"AA",x"4C",x"AA",x"4D",x"2D",x"D6",x"68",x"13",x"9B",x"31",x"95",x"86",x"A3",x"CF",x"74",x"D7",x"54",x"1A",x"B5",x"B1",x"E0",x"3D",x"13",x"6E",x"33",x"C6",x"0E",x"EB",x"42",x"B9",x"CD",x"98",x"1A",x"EC",x"2B",x"A3",x"36",x"63",x"2E",x"64",x"36",x"55",x"96",x"8E",x"B9",x"D0",x"D9",x"14",x"59",x"33",x"A6",x"42",x"67",x"4B",x"A4",x"C9",x"68",x"0A",x"99",x"4D",x"96",x"26",x"A3",x"2B",x"68",x"37",x"59",x"96",x"8C",x"BA",x"C1",x"D9",x"11",x"5A",x"D2",x"B2",x"0C",x"7F",x"54",x"BC",x"4E",x"4A",x"BC",x"FE",x"26",x"CA",x"26",x"29",x"F6",x"E2",x"93",x"A9",x"6A",x"97",x"B4",x"83",x"AA",x"36",x"13",x"53",x"CA",x"46",x"33",x"A2",x"33",x"4A",x"AA",x"1B",x"AE",x"88",x"AC",x"30",x"0C",x"E8",x"A0",x"C3",x"34",x"41",x"8F",x"57",x"28",x"6D",x"D3",x"3A",x"55",x"3E",x"6A",x"92",x"43",x"9B",x"94",x"4A",x"72",x"D6",x"1E",x"CD",x"D0",x"E1",x"E4",x"D6",x"79",x"D4",x"D3",x"4D",x"A2",x"5A",x"9B",x"51",x"CF",x"30",x"81",x"6C",x"6B",x"47",x"B5",x"7C",x"27",x"21",x"AF",x"1D",x"CD",x"F2",x"9B",x"88",x"D2",x"55",x"0D",x"5D",x"87",x"B1",x"59",x"EA",x"39",x"8C",x"66",x"E4",x"09",x"64",x"71",x"37",x"EA",x"15",x"2B",x"11",x"A5",x"EF",x"A8",x"77",x"CC",x"44",x"E4",x"2D",x"A5",x"D9",x"AE",x"1C",x"50",x"D7",x"A8",x"BA",x"B9",x"40",x"B4",x"4A",x"3D",x"92",x"A9",x"4A",x"91",x"A2",x"F5",x"88",x"17",x"0E",x"E3",x"F0",x"4D",x"23",x"69",x"2C",x"D4",x"DD",x"D7",x"B4",x"EA",x"98",x"70",x"13",x"75",x"AA",x"80",x"6B",x"D4",x"04",x"70",x"83",x"1A",x"01",x"1A",x"61",x"13",x"40",x"36",x"42",x"25",x"69",x"B9",x"54",x"2C",x"9C",x"B5",x"20",x"17",x"55",x"77",x"73",x"D6",x"BC",x"10",x"82",x"33",x"C5",x"59",x"73",x"A2",x"53",x"AF",x"46",x"AF",x"CD",x"4A",x"A2",x"87",x"53",x"3C",x"37",x"33",x"CA",x"1D",x"0D",x"4B",x"DD",x"AC",x"24",x"BB",x"22",x"B9",x"73",x"73",x"93",x"9C",x"92",x"F0",x"D6",x"2D",x"88",x"66",x"CA",x"D2",x"16",x"8D",x"AC",x"AA",x"36",x"0D",x"DB",x"3C",x"F2",x"21",x"DB",x"38",x"6D",x"CB",x"A8",x"BB",x"6F",x"16",x"F7",x"35",x"A3",x"EB",x"BE",x"94",x"3D",x"1B",x"8F",x"BE",x"87",x"32",x"8A",x"A8",x"3D",x"86",x"16",x"D3",x"28",x"BD",x"CA",x"18",x"BB",x"4D",x"15",x"F7",x"AA",x"6D",x"EC",x"B6",x"55",x"C2",x"B7",x"94",x"A9",x"DB",x"11",x"0E",x"DF",x"02",x"62",x"1D",x"B6",x"03",x"44",x"D6",x"20",x"20",x"59",x"B6",x"07",x"FF",
		x"60",x"02",x"A8",x"D3",x"5D",x"00",x"29",x"6A",x"10",x"20",x"64",x"49",x"17",x"C5",x"4C",x"95",x"21",x"2D",x"5B",x"94",x"AB",x"94",x"B9",x"CD",x"59",x"61",x"8D",x"65",x"9E",x"BA",x"66",x"45",x"35",x"A7",x"45",x"F8",x"D2",x"15",x"95",x"5C",x"16",x"E1",x"73",x"5B",x"9C",x"6B",x"58",x"44",x"CE",x"2D",x"71",x"AA",x"16",x"61",x"35",x"8F",x"00",x"BE",x"70",x"31",x"A0",x"14",x"CD",x"10",x"D6",x"D4",x"66",x"65",x"6B",x"52",x"D4",x"FC",x"B8",x"A5",x"2E",x"15",x"40",x"F5",x"E3",x"02",x"C8",x"6E",x"45",x"00",x"8B",x"5B",x"30",x"E0",x"5A",x"55",x"04",x"64",x"A4",x"AD",x"AA",x"C4",x"4C",x"AD",x"DD",x"89",x"C9",x"A3",x"08",x"F6",x"F4",x"D4",x"25",x"CD",x"95",x"D5",x"AD",x"EA",x"B4",x"A4",x"16",x"13",x"CD",x"9A",x"3B",x"92",x"9E",x"93",x"A9",x"6B",x"EE",x"48",x"BB",x"0B",x"A2",x"AE",x"A5",x"2D",x"1B",x"2D",x"89",x"CC",x"97",x"01",x"03",x"A2",x"17",x"13",x"40",x"0C",x"EC",x"A5",x"6A",x"D1",x"84",x"AB",x"AA",x"A4",x"B6",x"C7",x"40",x"AA",x"9A",x"92",x"EA",x"A2",x"84",x"EB",x"22",x"74",x"CA",x"03",x"EB",x"9C",x"06",x"AB",x"25",x"8F",x"F4",x"26",x"1D",x"6B",x"B7",x"2C",x"D1",x"1B",x"37",x"AE",x"53",x"D2",x"A8",x"AF",x"5D",x"78",x"6E",x"4B",x"93",x"B8",x"4E",x"E5",x"26",x"2D",x"4D",x"FC",x"26",x"94",x"1B",x"B7",x"34",x"CA",x"EB",x"14",x"5E",x"DC",x"D2",x"A8",x"AE",x"93",x"64",x"71",x"49",x"BC",x"BD",x"32",x"8A",x"C5",x"25",x"F1",x"E1",x"53",x"25",x"9B",x"96",x"D8",x"BB",x"2F",x"15",x"AF",x"53",x"22",x"EF",x"3E",x"58",x"A3",x"6E",x"89",x"A3",x"98",x"71",x"D2",x"B9",x"02",x"28",x"64",x"5A",x"00",x"85",x"CE",x"30",x"20",x"C9",x"6D",x"02",x"78",x"FB",x"85",x"00",x"6F",x"AF",x"4B",x"34",x"54",x"98",x"7A",x"36",x"6A",x"49",x"B5",x"2E",x"EC",x"F9",x"74",x"24",x"CD",x"8A",x"A9",x"F6",x"D2",x"92",x"4D",x"93",x"E2",x"A4",x"8D",x"04",x"B0",x"B8",x"B3",x"00",x"96",x"4A",x"4B",x"E1",x"60",x"E1",x"A2",x"DE",x"78",x"44",x"C5",x"B8",x"AA",x"D5",x"1C",x"13",x"17",x"27",x"26",x"B9",x"75",x"41",x"00",x"2D",x"3B",x"33",x"A0",x"87",x"94",x"14",x"EC",x"58",x"26",x"46",x"73",x"9B",x"BF",x"42",x"29",x"A9",x"2F",x"6D",x"C1",x"F4",x"AD",x"20",x"B9",x"B6",x"85",x"3D",x"26",x"41",x"64",x"DB",x"16",x"B7",x"18",x"84",x"E5",x"6D",x"5B",x"56",x"A3",x"13",x"8F",x"6E",x"6D",x"55",x"AD",x"4E",x"5A",x"BC",x"B9",x"75",x"35",x"25",x"73",x"73",x"9E",x"36",x"D5",x"12",x"AC",x"25",x"59",x"DB",x"9C",x"8B",x"B3",x"95",x"76",x"6D",x"6B",x"19",x"A1",x"1A",x"D4",x"A6",x"6C",x"65",x"9A",x"5A",x"50",x"DB",x"B4",x"E7",x"2E",x"62",x"2E",x"6B",x"C2",x"56",x"A6",x"5B",x"38",x"76",x"36",x"5B",x"69",x"CE",x"56",x"DC",x"FB",x"01",x"FF",
		x"60",x"4D",x"AE",x"BE",x"13",x"BB",x"93",x"0C",x"B1",x"9B",x"2E",x"B6",x"6D",x"3D",x"F8",x"AE",x"AB",x"C4",x"27",x"CE",x"E0",x"86",x"AE",x"51",x"CD",x"24",x"83",x"1D",x"A6",x"57",x"39",x"9D",x"0C",x"66",x"E8",x"5E",x"92",x"6C",x"32",x"98",x"A1",x"67",x"50",x"33",x"E9",x"60",x"86",x"EE",x"41",x"AD",x"24",x"83",x"19",x"AA",x"1A",x"B2",x"92",x"0C",x"66",x"C8",x"6A",x"AC",x"4C",x"3C",x"98",x"21",x"B3",x"B0",x"B3",x"F1",x"A0",x"07",x"CB",x"E6",x"CA",x"D4",x"83",x"6E",x"B4",x"4B",x"B2",x"DA",x"34",x"BA",x"B2",x"49",x"AE",x"DA",x"D2",x"E8",x"C2",x"36",x"B9",x"7A",x"F3",x"A0",x"2B",x"EB",x"A6",x"CE",x"35",x"83",x"CE",x"72",x"83",x"B3",x"D7",x"0C",x"26",x"8B",x"75",x"E9",x"5A",x"DA",x"98",x"C2",x"36",x"B8",x"6A",x"6D",x"63",x"0A",x"DD",x"E4",x"AA",x"B5",x"83",x"AD",x"64",x"8A",x"BA",x"1A",x"0F",x"B6",x"D1",x"2A",x"AA",x"6C",x"3D",x"B8",x"C6",x"3A",x"39",x"AA",x"F5",x"E0",x"1A",x"EB",x"E4",x"A8",x"C6",x"83",x"AF",x"6C",x"92",x"32",x"6B",x"37",x"BE",x"88",x"09",x"EA",x"AA",x"D3",x"F8",x"2C",x"26",x"A8",x"AB",x"4E",x"E3",x"33",x"9B",x"A2",x"A9",x"DA",x"4D",x"A8",x"B8",x"1A",x"A7",x"1B",x"35",x"A1",x"E1",x"18",x"9C",x"69",x"D5",x"C4",x"42",x"AB",x"B1",x"A7",x"71",x"93",x"B2",x"1C",x"C7",x"9A",x"C6",x"45",x"CA",x"72",x"03",x"66",x"6A",x"17",x"B9",x"88",x"49",x"D8",x"49",x"52",x"E4",x"AC",x"D6",x"A1",x"B6",x"49",x"51",x"B2",x"3E",x"83",x"DC",x"C6",x"45",x"2D",x"62",x"0A",x"7A",x"92",x"24",x"B5",x"F0",x"29",x"88",x"49",x"93",x"B4",x"2C",x"27",x"C1",x"D7",x"6D",x"D2",x"B3",x"DA",x"80",x"A8",x"A4",x"C1",x"2C",x"74",x"1A",x"A3",x"EC",x"04",x"AB",x"91",x"5C",x"88",x"76",x"1C",x"EC",x"42",x"6A",x"C0",x"C7",x"49",x"B0",x"2B",x"EE",x"21",x"ED",x"38",x"C1",x"E9",x"C8",x"96",x"B4",x"ED",x"04",x"B7",x"E0",x"1E",x"B2",x"8E",x"E3",x"BC",x"44",x"B7",x"31",x"26",x"8E",x"F3",x"13",x"9D",x"C1",x"98",x"A4",x"21",x"A8",x"B4",x"86",x"24",x"9A",x"88",x"20",x"F1",x"1E",x"72",x"9F",x"FA",x"00",x"FF",
		x"60",x"43",x"19",x"7C",x"02",x"7B",x"93",x"0D",x"79",x"D1",x"2C",x"AE",x"49",x"3A",x"A4",x"C5",x"B3",x"38",x"26",x"EE",x"90",x"96",x"E8",x"A2",x"18",x"BB",x"43",x"EA",x"72",x"1D",x"BB",x"DD",x"0C",x"A9",x"E9",x"31",x"DA",x"F0",x"34",x"A4",x"AA",x"DB",x"78",x"DD",x"F5",x"90",x"9B",x"1C",x"E3",x"0D",x"27",x"43",x"69",x"BC",x"83",x"36",x"93",x"0E",x"B5",x"C8",x"31",x"BD",x"72",x"3B",x"D4",x"2C",x"C7",x"EC",x"33",x"ED",x"D0",x"0A",x"9F",x"90",x"EF",x"A4",x"43",x"CF",x"62",x"4C",x"BF",x"9D",x"0C",x"BD",x"C8",x"51",x"FE",x"4D",x"3A",x"8D",x"61",x"17",x"B9",x"4A",x"3B",x"6E",x"87",x"53",x"F9",x"1A",x"6D",x"3B",x"1D",x"4E",x"27",x"9D",x"38",x"E3",x"74",x"B8",x"8D",x"4E",x"E0",x"B6",x"93",x"E1",x"36",x"36",x"8E",x"33",x"4E",x"86",x"D7",x"D8",x"04",x"CE",x"B8",x"1E",x"7E",x"C7",x"DD",x"34",x"ED",x"66",x"F8",x"15",x"4F",x"EA",x"B6",x"E3",x"11",x"54",x"36",x"4E",x"B7",x"4E",x"46",x"58",x"E9",x"38",x"DD",x"26",x"1D",x"51",x"25",x"13",x"B4",x"9B",x"74",x"44",x"8D",x"76",x"C2",x"6E",x"D2",x"91",x"0C",x"36",x"05",x"31",x"4D",x"47",x"F6",x"A4",x"B6",x"72",x"D5",x"19",x"F9",x"15",x"39",x"82",x"51",x"77",x"E4",x"57",x"C4",x"38",x"C4",x"DC",x"51",x"5C",x"65",x"1D",x"90",x"73",x"47",x"79",x"94",x"8F",x"63",x"36",x"19",x"D5",x"91",x"BE",x"0A",x"DD",x"74",x"54",x"47",x"E9",x"18",x"54",x"93",x"51",x"5D",x"65",x"63",x"D0",x"4D",x"46",x"75",x"95",x"8E",x"41",x"37",x"19",x"F5",x"33",x"D2",x"09",x"D5",x"64",x"D4",x"CF",x"C8",x"04",x"56",x"E3",x"D1",x"3C",x"23",x"13",x"98",x"4D",x"47",x"F3",x"8C",x"8C",x"63",x"2E",x"69",x"ED",x"93",x"3C",x"41",x"D5",x"64",x"B4",x"4F",x"C9",x"04",x"64",x"D3",x"D1",x"3C",x"A9",x"E3",x"58",x"4D",x"46",x"73",x"99",x"8F",x"E2",x"D4",x"69",x"CD",x"21",x"3E",x"82",x"53",x"A7",x"35",x"1B",x"E7",x"30",x"6D",x"9D",x"56",x"6F",x"14",x"A3",x"BC",x"71",x"5A",x"D5",x"E0",x"8C",x"F8",x"DA",x"49",x"55",x"92",x"27",x"B2",x"AD",x"24",x"D5",x"95",x"4E",x"C2",x"94",x"E3",x"D4",x"74",x"D2",x"89",x"D9",x"8A",x"5D",x"DB",x"D8",x"14",x"66",x"29",x"7E",x"FF",
		x"60",x"83",x"3E",x"CA",x"D3",x"82",x"D8",x"0C",x"7A",x"99",x"54",x"2B",x"52",x"3A",x"98",x"65",x"9D",x"75",x"DC",x"CD",x"60",x"A7",x"33",x"B5",x"61",x"25",x"83",x"1D",x"42",x"2D",x"47",x"DC",x"0E",x"76",x"68",x"B5",x"6C",x"74",x"3B",x"98",x"25",x"CD",x"A2",x"59",x"CD",x"60",x"B6",x"72",x"89",x"11",x"37",x"83",x"DD",x"C2",x"2D",x"5A",x"95",x"0C",x"EE",x"48",x"F7",x"58",x"52",x"32",x"B8",x"C5",x"DC",x"A3",x"C5",x"EE",x"E0",x"27",x"8B",x"C8",x"C2",x"A4",x"43",x"98",x"34",x"33",x"13",x"D3",x"0D",x"61",x"92",x"CC",x"08",x"4C",x"37",x"84",x"49",x"A2",x"22",x"29",x"ED",x"10",x"1B",x"EB",x"8E",x"80",x"B6",x"43",x"AA",x"7C",x"BA",x"1C",x"BA",x"0C",x"A9",x"F1",x"AC",x"4A",x"E8",x"32",x"E4",x"8A",x"32",x"AB",x"39",x"CD",x"50",x"0A",x"AA",x"CE",x"E2",x"B4",x"43",x"2D",x"38",x"72",x"46",x"5C",x"0F",x"B5",x"12",x"F3",x"5D",x"49",x"3C",x"F4",x"C9",x"C4",x"7D",x"C5",x"F1",x"30",x"3A",x"8D",x"8A",x"A4",x"34",x"C3",x"6C",x"BC",x"3B",x"02",x"D2",x"0C",x"A3",x"F3",x"EA",x"08",x"48",x"3B",x"CC",x"C6",x"7B",x"B2",x"C0",x"E9",x"B0",x"AB",x"A8",x"CA",x"80",x"A6",x"C3",x"CD",x"A2",x"2B",x"1D",x"DB",x"0C",x"B7",x"D1",x"AC",x"28",x"6C",x"3B",x"DC",x"4A",x"B3",x"B2",x"38",x"DD",x"F0",x"0A",x"CD",x"CA",x"A2",x"B6",x"C3",x"AB",x"D4",x"B3",x"07",x"BB",x"0E",x"BF",x"08",x"CF",x"0A",x"EC",x"3A",x"FC",x"CC",x"BB",x"CC",x"A9",x"DF",x"F0",x"93",x"EC",x"32",x"E3",x"75",x"C3",x"4F",x"2C",x"6A",x"86",x"D3",x"8E",x"20",x"B1",x"A8",x"59",x"4E",x"3A",x"82",x"C8",x"B2",x"67",x"39",x"E9",x"08",x"33",x"89",x"EA",x"E5",x"D4",x"23",x"2A",x"D4",x"B2",x"97",x"DD",x"8C",x"A8",x"62",x"EB",x"1A",x"76",x"32",x"A2",x"46",x"AC",x"6A",x"D9",x"C9",x"88",x"1B",x"B3",x"AC",x"46",x"2F",x"23",x"6E",x"CC",x"2B",x"12",x"B2",x"8E",x"A4",x"51",x"6F",x"0F",x"F2",x"3A",x"92",x"46",x"BD",x"23",x"C9",x"CB",x"48",x"1A",x"8D",x"CE",x"C4",x"2C",x"23",x"ED",x"C4",x"3B",x"83",x"B5",x"8C",x"B4",x"91",x"98",x"08",x"F2",x"3A",x"B2",x"86",x"A3",x"D3",x"D9",x"EB",x"C8",x"3A",x"F6",x"AA",x"14",x"BE",x"23",x"EB",x"C4",x"AA",x"5A",x"B4",x"8C",x"6C",x"60",x"ED",x"4E",x"E5",x"32",x"B2",x"8E",x"B5",x"7A",x"54",x"CD",x"C8",x"3A",x"D6",x"EC",x"51",x"36",x"23",x"1B",x"D0",x"6A",x"DA",x"D8",x"8C",x"BC",x"43",x"CF",x"69",x"E5",x"3A",x"F2",x"8E",x"3C",x"A7",x"95",x"EB",x"C8",x"3B",x"B6",x"98",x"51",x"AE",x"23",x"EF",x"30",x"6A",x"4A",x"B9",x"8E",x"A2",x"C2",x"EC",x"4E",x"D1",x"3A",x"8A",x"06",x"B2",x"26",x"54",x"EF",x"2A",x"0A",x"9A",x"72",x"B1",x"BC",x"A3",x"AC",x"70",x"DB",x"28",x"F2",x"8D",x"32",x"A3",x"AD",x"10",x"CD",x"3B",x"CA",x"0A",x"AF",x"9C",x"2D",x"EF",x"A8",x"2A",x"9C",x"6C",x"11",x"BF",x"A3",x"6E",x"24",x"73",x"9C",x"35",x"A7",x"36",x"A9",x"C9",x"26",x"4E",x"E3",x"DA",x"46",x"22",x"DA",x"C8",x"31",x"02",x"02",x"3D",x"47",x"40",x"E0",x"1B",x"08",x"88",x"7C",x"02",x"01",x"99",x"A5",x"3F",x"FF",
		x"60",x"8D",x"CD",x"D6",x"BD",x"52",x"D7",x"0C",x"A1",x"24",x"AD",x"30",x"6F",x"32",x"F8",x"12",x"32",x"DC",x"69",x"C9",x"60",x"8B",x"37",x"CF",x"E0",x"B5",x"83",x"2D",x"DE",x"AC",x"8A",x"D6",x"0D",x"AE",x"3A",x"F1",x"2A",x"5E",x"3D",x"F8",x"12",x"3D",x"32",x"71",x"4D",x"11",x"73",x"B4",x"8C",x"E0",x"35",x"43",x"2A",x"51",x"33",x"83",x"96",x"0C",x"B9",x"06",x"8B",x"4C",x"6C",x"3B",x"94",x"1A",x"2D",x"2B",x"B1",x"E9",x"50",x"4B",x"D2",x"4A",x"E7",x"35",x"4D",x"CB",x"49",x"3B",x"5C",x"56",x"37",x"35",x"47",x"AD",x"74",x"5E",x"DC",x"D4",x"12",x"35",x"B3",x"70",x"CD",x"D0",x"8A",x"B3",x"8C",x"A6",x"B5",x"43",x"AB",x"D6",x"C2",x"87",x"D3",x"35",x"3D",x"39",x"CF",x"28",x"69",x"57",x"F4",x"E8",x"A2",x"A2",x"3C",x"69",x"D1",x"93",x"CB",x"B4",x"F2",x"A4",x"45",x"CF",x"21",x"C2",x"5D",x"DA",x"15",x"23",x"F9",x"70",x"4F",x"6B",x"9B",x"F4",x"12",x"34",x"C3",x"A5",x"49",x"32",x"93",x"0B",x"D7",x"B0",x"A6",x"C9",x"48",x"C1",x"5D",x"C3",x"92",x"24",x"23",x"15",x"37",x"0D",x"6D",x"52",x"8C",x"14",x"C2",x"35",x"AC",x"4D",x"32",x"52",x"4C",x"D3",x"B0",x"C6",x"C1",x"4A",x"2E",x"42",x"C2",x"53",x"3B",x"3B",x"EB",x"08",x"0D",x"4B",x"EA",x"EC",x"62",x"D5",x"C3",x"38",x"8D",x"71",x"8B",x"56",x"CF",x"14",x"39",x"0F",x"FF",
		x"60",x"45",x"CA",x"5E",x"3D",x"A3",x"63",x"0F",x"A1",x"5A",x"F5",x"F2",x"88",x"35",x"F8",x"6A",x"5D",x"53",x"A3",x"D6",x"60",x"9A",x"2B",x"77",x"D1",x"AD",x"83",x"EE",x"BE",x"23",x"85",x"B7",x"0C",x"A6",x"B9",x"B4",x"50",x"5B",x"33",x"F8",x"EC",x"D5",x"3C",x"6A",x"F4",x"E0",x"6B",x"D0",x"50",x"EB",x"D9",x"43",x"28",x"5E",x"CD",x"AD",x"97",x"0C",x"31",x"7B",x"53",x"B7",x"5E",x"37",x"E4",x"EA",x"C4",x"43",x"7A",x"EE",x"50",x"8A",x"35",x"0D",x"AB",x"25",x"43",x"29",x"D6",x"34",x"BC",x"E6",x"0C",x"AD",x"78",x"35",x"B5",x"9A",x"3D",x"B4",x"6C",x"55",x"DD",x"63",x"76",x"D3",x"B2",x"36",x"F3",x"8C",x"DB",x"4D",x"CF",x"46",x"DC",x"2D",x"6E",x"17",x"BD",x"58",x"4E",x"D7",x"BA",x"5C",x"F4",x"6C",x"39",x"5D",x"F3",x"72",x"35",x"9A",x"99",x"83",x"AA",x"5A",x"CE",x"2E",x"56",x"0A",x"EA",x"AA",x"39",x"25",x"D9",x"D9",x"71",x"AA",x"D4",x"94",x"E4",x"26",x"19",x"AA",x"65",x"B3",x"83",x"1B",x"AD",x"A9",x"45",x"D4",x"74",x"7E",x"B6",x"AA",x"2E",x"BE",x"D0",x"04",x"D5",x"88",x"A9",x"F3",x"42",x"13",x"55",x"65",x"2A",x"A1",x"29",x"59",x"52",x"7D",x"28",x"09",x"B6",x"7A",x"FF",
		x"60",x"83",x"5B",x"9E",x"4B",x"5D",x"88",x"0D",x"6E",x"5A",x"4D",x"2E",x"15",x"37",x"F8",x"E5",x"D5",x"31",x"23",x"EC",x"10",x"BA",x"16",x"93",x"71",x"6B",x"43",x"EC",x"8A",x"5D",x"27",x"AC",x"0D",x"B1",x"0B",x"0A",x"9F",x"8C",x"36",x"C4",x"EE",x"D4",x"6D",x"54",x"EC",x"10",x"A6",x"61",x"97",x"0E",x"63",x"43",x"98",x"56",x"9C",x"27",x"CC",x"0D",x"61",x"59",x"71",x"1E",x"37",x"3B",x"A4",x"65",x"39",x"65",x"4D",x"EC",x"90",x"96",x"E1",x"D4",x"76",x"B3",x"43",x"9E",x"9A",x"52",x"D7",x"A4",x"0E",x"65",x"08",x"69",x"1D",x"96",x"3F",x"94",x"21",x"A5",x"AD",x"59",x"FA",x"50",x"87",x"90",x"B6",x"66",x"F9",x"43",x"1B",x"82",x"DB",x"5A",x"A4",x"0F",x"BD",x"0B",x"1D",x"6B",x"A2",x"3F",x"8C",x"26",x"6C",x"AC",x"89",x"FE",x"30",x"AA",x"B0",x"B1",x"26",x"FA",x"C3",x"6C",x"42",x"DB",x"86",x"E8",x"0F",x"AB",x"71",x"49",x"5B",x"95",x"3F",x"9C",x"C6",x"39",x"F4",x"42",x"DA",x"70",x"BB",x"E0",x"B6",x"51",x"69",x"C3",x"6B",x"42",x"DB",x"86",x"E5",x"0F",x"B7",x"09",x"1B",x"6B",x"92",x"3F",x"BC",x"2A",x"6C",x"AC",x"50",x"FE",x"F0",x"8A",x"F4",x"B5",x"46",x"79",x"CD",x"CF",x"D2",x"C7",x"1A",x"95",x"B5",x"20",x"4B",x"6B",x"1F",x"52",x"D6",x"C2",x"C2",x"6D",x"AC",x"59",x"79",x"0B",x"2B",x"97",x"B1",x"65",x"7B",x"2D",x"2C",x"DC",x"C6",x"47",x"9C",x"B5",x"B0",x"70",x"1D",x"5F",x"51",x"DE",x"A2",x"2C",x"B4",x"FD",x"44",x"79",x"8B",x"B2",x"D4",x"8A",x"61",x"E5",x"23",x"CA",x"C2",x"C7",x"92",x"95",x"B7",x"38",x"0B",x"1F",x"2B",x"72",x"DE",x"E2",x"24",x"6C",x"7C",x"C8",x"7D",x"8B",x"13",x"D7",x"CE",x"0F",x"69",x"2D",x"4D",x"4C",x"3B",x"2F",x"A4",x"B5",x"34",x"33",x"E9",x"D8",x"14",x"D7",x"D2",x"CC",x"A4",x"E3",x"5C",x"5A",x"4B",x"0B",x"E3",x"F1",x"75",x"71",x"2D",x"AB",x"9C",x"DB",x"C7",x"C4",x"B5",x"BC",x"0A",x"29",x"6F",x"95",x"DE",x"F2",x"2A",x"64",x"AC",x"59",x"7E",x"CB",x"1B",x"E7",x"F1",x"54",x"E9",x"2D",x"AF",x"42",x"C6",x"4B",x"A4",x"B7",x"A2",x"70",x"69",x"1F",x"56",x"DE",x"8A",x"CA",x"B9",x"A3",x"54",x"7A",x"2B",x"2B",x"E7",x"C9",x"54",x"E9",x"AD",x"AC",x"5C",x"26",x"43",x"A4",x"B7",x"B2",x"31",x"E9",x"4A",x"11",x"DF",x"AA",x"C6",x"B8",x"B2",x"5D",x"78",x"AB",x"1A",x"E7",x"CA",x"09",x"E3",x"AD",x"EA",x"9C",x"AA",x"DA",x"8D",x"B5",x"AA",x"73",x"CA",x"9A",x"30",x"D6",x"AA",x"CE",x"38",x"6B",x"C2",x"58",x"AB",x"3A",x"E5",x"AA",x"71",x"63",x"AD",x"EE",x"94",x"B3",x"26",x"82",x"B5",x"BA",x"53",x"CE",x"DC",x"30",x"D6",x"EA",x"46",x"39",x"73",x"C3",x"58",x"AB",x"3B",x"E3",x"C8",x"C9",x"60",x"AD",x"6E",x"44",x"AA",x"26",x"8C",x"B5",x"A6",x"62",x"E9",x"1E",x"33",x"DE",x"EA",x"8A",x"A5",x"6B",x"CC",x"78",x"6B",x"2B",x"D6",x"CE",x"56",x"F3",x"AD",x"2D",x"C8",x"27",x"9C",x"E2",x"F7",x"B6",x"B5",x"05",x"C5",x"44",x"50",x"FC",x"D6",x"56",x"68",x"93",x"41",x"D1",x"5B",x"17",x"59",x"8D",x"07",x"25",x"6F",x"7D",x"C3",x"52",x"D5",x"6A",x"BC",x"0C",x"59",x"64",x"57",x"B0",x"F4",x"30",x"24",x"95",x"95",x"85",x"F2",x"D4",x"D4",x"A8",x"96",x"0F",x"49",x"7B",x"FF",
		x"60",x"4D",x"AE",x"BE",x"13",x"BB",x"93",x"0C",x"B1",x"9B",x"2E",x"B6",x"6D",x"3D",x"F8",x"AE",x"AB",x"C4",x"27",x"CE",x"E0",x"86",x"AE",x"51",x"CD",x"24",x"83",x"1D",x"A6",x"57",x"39",x"9D",x"0C",x"66",x"E8",x"5E",x"92",x"6C",x"32",x"98",x"A1",x"67",x"50",x"33",x"E9",x"60",x"86",x"EE",x"41",x"AD",x"24",x"83",x"19",x"AA",x"1A",x"B2",x"92",x"0C",x"66",x"C8",x"6A",x"AC",x"4C",x"3C",x"98",x"21",x"B3",x"B0",x"B3",x"F1",x"A0",x"07",x"CB",x"E6",x"CA",x"D4",x"83",x"6E",x"B4",x"4B",x"B2",x"DA",x"34",x"BA",x"B2",x"49",x"AE",x"DA",x"D2",x"E8",x"C2",x"36",x"B9",x"7A",x"F3",x"A0",x"2B",x"EB",x"A6",x"CE",x"35",x"83",x"CE",x"72",x"83",x"B3",x"D7",x"0C",x"26",x"8B",x"75",x"E9",x"5A",x"DA",x"98",x"C2",x"36",x"B8",x"6A",x"6D",x"63",x"0A",x"DD",x"E4",x"AA",x"B5",x"83",x"AD",x"64",x"8A",x"BA",x"1A",x"0F",x"B6",x"D1",x"2A",x"AA",x"6C",x"3D",x"B8",x"C6",x"3A",x"39",x"AA",x"F5",x"E0",x"1A",x"EB",x"E4",x"A8",x"C6",x"83",x"AF",x"6C",x"92",x"32",x"6B",x"37",x"BE",x"88",x"09",x"EA",x"AA",x"D3",x"F8",x"2C",x"26",x"A8",x"AB",x"4E",x"E3",x"33",x"9B",x"A2",x"A9",x"DA",x"4D",x"A8",x"B8",x"1A",x"A7",x"1B",x"35",x"A1",x"E1",x"18",x"9C",x"69",x"D5",x"C4",x"42",x"AB",x"B1",x"A7",x"71",x"93",x"B2",x"1C",x"C7",x"9A",x"C6",x"45",x"CA",x"72",x"03",x"66",x"6A",x"17",x"B9",x"88",x"49",x"D8",x"49",x"52",x"E4",x"AC",x"D6",x"A1",x"B6",x"49",x"51",x"B2",x"3E",x"83",x"DC",x"C6",x"45",x"2D",x"62",x"0A",x"7A",x"92",x"24",x"B5",x"F0",x"29",x"88",x"49",x"93",x"B4",x"2C",x"27",x"C1",x"D7",x"6D",x"D2",x"B3",x"DA",x"80",x"A8",x"A4",x"C1",x"2C",x"74",x"1A",x"A3",x"EC",x"04",x"AB",x"91",x"5C",x"88",x"76",x"1C",x"EC",x"42",x"6A",x"C0",x"C7",x"49",x"B0",x"2B",x"EE",x"21",x"ED",x"38",x"C1",x"E9",x"C8",x"96",x"B4",x"ED",x"04",x"B7",x"E0",x"1E",x"B2",x"8E",x"E3",x"BC",x"44",x"B7",x"31",x"26",x"8E",x"F3",x"13",x"9D",x"C1",x"98",x"A4",x"21",x"A8",x"B4",x"86",x"24",x"9A",x"88",x"20",x"F1",x"1E",x"72",x"9F",x"FA",x"00",x"FF",
		x"60",x"43",x"19",x"7C",x"02",x"7B",x"93",x"0D",x"79",x"D1",x"2C",x"AE",x"49",x"3A",x"A4",x"C5",x"B3",x"38",x"26",x"EE",x"90",x"96",x"E8",x"A2",x"18",x"BB",x"43",x"EA",x"72",x"1D",x"BB",x"DD",x"0C",x"A9",x"E9",x"31",x"DA",x"F0",x"34",x"A4",x"AA",x"DB",x"78",x"DD",x"F5",x"90",x"9B",x"1C",x"E3",x"0D",x"27",x"43",x"69",x"BC",x"83",x"36",x"93",x"0E",x"B5",x"C8",x"31",x"BD",x"72",x"3B",x"D4",x"2C",x"C7",x"EC",x"33",x"ED",x"D0",x"0A",x"9F",x"90",x"EF",x"A4",x"43",x"CF",x"62",x"4C",x"BF",x"9D",x"0C",x"BD",x"C8",x"51",x"FE",x"4D",x"3A",x"8D",x"61",x"17",x"B9",x"4A",x"3B",x"6E",x"87",x"53",x"F9",x"1A",x"6D",x"3B",x"1D",x"4E",x"27",x"9D",x"38",x"E3",x"74",x"B8",x"8D",x"4E",x"E0",x"B6",x"93",x"E1",x"36",x"36",x"8E",x"33",x"4E",x"86",x"D7",x"D8",x"04",x"CE",x"B8",x"1E",x"7E",x"C7",x"DD",x"34",x"ED",x"66",x"F8",x"15",x"4F",x"EA",x"B6",x"E3",x"11",x"54",x"36",x"4E",x"B7",x"4E",x"46",x"58",x"E9",x"38",x"DD",x"26",x"1D",x"51",x"25",x"13",x"B4",x"9B",x"74",x"44",x"8D",x"76",x"C2",x"6E",x"D2",x"91",x"0C",x"36",x"05",x"31",x"4D",x"47",x"F6",x"A4",x"B6",x"72",x"D5",x"19",x"F9",x"15",x"39",x"82",x"51",x"77",x"E4",x"57",x"C4",x"38",x"C4",x"DC",x"51",x"5C",x"65",x"1D",x"90",x"73",x"47",x"79",x"94",x"8F",x"63",x"36",x"19",x"D5",x"91",x"BE",x"0A",x"DD",x"74",x"54",x"47",x"E9",x"18",x"54",x"93",x"51",x"5D",x"65",x"63",x"D0",x"4D",x"46",x"75",x"95",x"8E",x"41",x"37",x"19",x"F5",x"33",x"D2",x"09",x"D5",x"64",x"D4",x"CF",x"C8",x"04",x"56",x"E3",x"D1",x"3C",x"23",x"13",x"98",x"4D",x"47",x"F3",x"8C",x"8C",x"63",x"2E",x"69",x"ED",x"93",x"3C",x"41",x"D5",x"64",x"B4",x"4F",x"C9",x"04",x"64",x"D3",x"D1",x"3C",x"A9",x"E3",x"58",x"4D",x"46",x"73",x"99",x"8F",x"E2",x"D4",x"69",x"CD",x"21",x"3E",x"82",x"53",x"A7",x"35",x"1B",x"E7",x"30",x"6D",x"9D",x"56",x"6F",x"14",x"A3",x"BC",x"71",x"5A",x"D5",x"E0",x"8C",x"F8",x"DA",x"49",x"55",x"92",x"27",x"B2",x"AD",x"24",x"D5",x"95",x"4E",x"C2",x"94",x"E3",x"D4",x"74",x"D2",x"89",x"D9",x"8A",x"5D",x"DB",x"D8",x"14",x"66",x"29",x"7E",x"FF"
	);

	-- Clock period for 640KHz
	constant CLK_period : time := 1 ms / 640;

begin
	uut: entity work.TMS5220 port map (
		I_OSC    => CLK,
		I_ENA    => '1',
		I_WSn    => I_WSn,
		I_RSn    => I_RSn,
		I_DATA   => I_DATA,
		I_TEST   => I_TEST,
		I_DBUS   => I_DBUS,
		O_DBUS   => O_DBUS,
		O_RDYn   => O_RDYn,
		O_INTn   => O_INTn,
		O_M0     => O_M0,
		O_M1     => O_M1,
		O_ADD8   => O_ADD8,
		O_ADD4   => O_ADD4,
		O_ADD2   => O_ADD2,
		O_ADD1   => O_ADD1,
		O_ROMCLK => O_ROMCLK,
		O_T11    => O_T11,
		O_IO     => O_IO,
		O_PRMOUT => O_PRMOUT,
		O_SPKR   => O_SPKR
	);

	-- Clock process definitions
	p_CLK : process
	begin
		CLK <= '0';
		wait for CLK_period/2;
		CLK <= '1';
		wait for CLK_period/2;
	end process;

	-- Stimulus process - state machine
	stim_proc: process
	begin
		wait until rising_edge(CLK);
		case state is
			when 0 =>				-- init signal levels
				I_DATA  <= '1';
				I_TEST  <= '1';
				index   <= 0;
				current <= 0;
				offset  <= 0;
				state   <= state + 1;

				I_WSn   <= '0';		-- chip reset
				I_RSn   <= '0';

			when 1 =>
				I_WSn   <= '1';		-- release reset
				I_RSn   <= '1';
				state   <= state + 1;

			-- read status
			when 2 =>				-- assert RSn
				I_RSn <= '0';
				state <= state + 1;

			when 3 =>
				I_RSn <= '1';		-- deassert RSn
				state <= state + 1;

			when 4 =>				-- if Talk Status
				if (O_DBUS(7) = '1') then
					state <= 8;
				else
					state <= state + 1;
				end if;

			when 5 =>				-- if Buffer Low
				if (index < SIZES(current)) and (O_DBUS(6) = '1') then
					I_DBUS <= DATA(offset + index);
					index  <= index + 1;
					state  <= state + 1;
				else
					state <= 2;
				end if;

			-- write data
			when 6 =>				-- assert WSn
				I_WSn  <= '0';
				state  <= state + 1;

			when 7 =>				-- deassert WSn
				I_WSn <= '1';
				state <= 2;

			-- read status
			when 8 =>				-- assert RSn
				I_RSn <= '0';
				state <= state + 1;

			when 9 =>
				I_RSn <= '1';		-- deassert RSn
				state <= state + 1;

			when 10 =>				-- if Talk Status
				if (O_DBUS(7) = '1') then
					state <= 12;
				else
					index   <= 0;
					offset  <= offset + index;
					current <= current + 1;
					state   <= state + 1;
				end if;

			when 11 =>				-- if more sounds
				if (current < MAXSOUNDS) then
					state   <= 2;
				end if;

			when 12 =>				-- if Buffer Low
				if (index < SIZES(current)) and (O_DBUS(6) = '1') then
					index  <= index + 1;
					I_DBUS <= DATA(offset + index);
					state   <= state + 1;
				else
					state <= 8;
				end if;

			-- write data
			when 13 =>				-- assert WSn
				I_WSn  <= '0';
				state  <= state + 1;

			when 14 =>				-- deassert WSn
				I_WSn <= '1';
				state <= 8;

			when others => null;	-- end state
		end case;
	end process;
end;
